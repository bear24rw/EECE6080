magic
tech scmos
timestamp 1383792416
<< metal1 >>
rect -1 162 3 165
rect -8 153 -1 156
rect -1 109 2343 113
<< m2contact >>
rect -5 161 -1 165
rect 10 117 14 121
rect -5 109 -1 113
rect 2343 109 2347 113
rect 10 1 14 5
<< metal2 >>
rect -5 113 -1 161
rect 10 121 14 128
rect 101 93 105 129
rect 257 93 261 129
rect 413 93 417 129
rect 569 93 573 129
rect 725 93 729 129
rect 881 93 885 129
rect 1037 93 1041 129
rect 1193 93 1197 129
rect 1349 93 1353 129
rect 1505 93 1509 129
rect 1661 93 1665 129
rect 1817 93 1821 129
rect 1973 93 1977 129
rect 2129 93 2133 129
rect 2285 93 2289 129
rect 2343 46 2347 109
rect 10 5 14 16
<< end >>
