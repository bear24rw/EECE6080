magic
tech scmos
timestamp 1383629942
<< metal1 >>
rect 31 37 39 40
<< m2contact >>
rect 11 46 15 50
use BUFX4  BUFX4_0
timestamp 1383629942
transform 1 0 9 0 1 3
box -9 -3 37 105
<< end >>
