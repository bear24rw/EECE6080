magic
tech scmos
timestamp 1383914834
<< metal1 >>
rect 1020 3982 1044 3991
rect 1053 3982 1311 3991
rect 1320 3982 1344 3991
rect 1353 3982 1857 3991
rect 1866 3982 2157 3991
rect 1620 3964 1911 3973
rect 1920 3964 2148 3973
rect 2139 3879 2148 3964
rect 2157 3899 2166 3982
rect 2302 3950 2398 4000
rect 2520 3982 2544 3991
rect 2553 3982 2811 3991
rect 2820 3982 2844 3991
rect 2853 3982 3111 3991
rect 3120 3982 3144 3991
rect 3153 3982 3411 3991
rect 3420 3982 3444 3991
rect 3453 3982 3957 3991
rect 2303 3949 2397 3950
rect 2304 3948 2396 3949
rect 2305 3947 2395 3948
rect 2306 3946 2394 3947
rect 2307 3945 2393 3946
rect 2308 3944 2392 3945
rect 2309 3943 2391 3944
rect 2310 3942 2390 3943
rect 2311 3941 2389 3942
rect 2312 3940 2388 3941
rect 2313 3939 2387 3940
rect 2314 3938 2386 3939
rect 2315 3937 2385 3938
rect 2316 3936 2384 3937
rect 2317 3935 2383 3936
rect 2318 3934 2382 3935
rect 2319 3933 2381 3934
rect 2320 3932 2380 3933
rect 2321 3931 2379 3932
rect 2322 3930 2378 3931
rect 2323 3929 2377 3930
rect 2324 3928 2376 3929
rect 2325 3927 2375 3928
rect 2326 3926 2374 3927
rect 2327 3925 2373 3926
rect 2328 3924 2372 3925
rect 2329 3923 2371 3924
rect 2330 3922 2370 3923
rect 2331 3921 2369 3922
rect 2332 3920 2368 3921
rect 2333 3919 2367 3920
rect 2334 3918 2366 3919
rect 2335 3917 2365 3918
rect 2336 3916 2364 3917
rect 2337 3915 2363 3916
rect 2338 3914 2362 3915
rect 2339 3913 2361 3914
rect 2340 3912 2360 3913
rect 2341 3911 2359 3912
rect 2342 3910 2358 3911
rect 2343 3909 2357 3910
rect 2344 3908 2356 3909
rect 2345 3879 2355 3908
rect 2511 3899 2520 3982
rect 3982 3973 3991 3980
rect 2529 3964 3711 3973
rect 3720 3964 3991 3973
rect 2529 3879 2538 3964
rect 1009 3420 1018 3711
rect 3982 3689 3991 3734
rect 3982 3656 3991 3680
rect 3982 3566 3991 3647
rect 3900 3556 3991 3566
rect 1018 3411 1101 3420
rect 3900 3380 3982 3389
rect 1018 3144 1101 3153
rect 1018 3057 1101 3066
rect 3900 2834 3982 2843
rect 1018 2811 1121 2820
rect 3880 2780 3982 2789
rect 3900 2534 3982 2543
rect 1018 2511 1101 2520
rect 3880 2480 3982 2489
rect 3900 2234 3982 2243
rect 1018 2211 1101 2220
rect 3880 2180 3982 2189
rect 3900 1934 3982 1943
rect 1018 1911 1101 1920
rect 3880 1880 3982 1889
rect 3900 1634 3982 1643
rect 1018 1611 1101 1620
rect 3880 1580 3982 1589
rect 3900 1334 3982 1343
rect 1018 1311 1101 1320
rect 1009 1053 1018 1311
rect 3880 1280 3982 1289
rect 2439 1036 2448 1121
rect 1026 1027 1311 1036
rect 1320 1027 1611 1036
rect 1620 1027 1911 1036
rect 1920 1027 2211 1036
rect 2220 1027 2448 1036
rect 1026 1018 1035 1027
rect 2457 1018 2466 1141
rect 1266 1009 1557 1018
rect 1566 1009 1857 1018
rect 1866 1009 2157 1018
rect 2166 1009 2457 1018
rect 2793 1018 2802 1141
rect 2811 1036 2820 1121
rect 2820 1027 3111 1036
rect 3120 1027 3411 1036
rect 3420 1027 3711 1036
rect 3982 1018 3991 1034
rect 2793 1009 3057 1018
rect 3066 1009 3357 1018
rect 3366 1009 3657 1018
rect 3666 1009 3957 1018
rect 3966 1009 3991 1018
<< m2contact >>
rect 1011 3982 1020 3991
rect 1044 3982 1053 3991
rect 1311 3982 1320 3991
rect 1344 3982 1353 3991
rect 1857 3982 1866 3991
rect 2157 3982 2166 3991
rect 1611 3964 1620 3973
rect 1911 3964 1920 3973
rect 2511 3982 2520 3991
rect 2544 3982 2553 3991
rect 2811 3982 2820 3991
rect 2844 3982 2853 3991
rect 3111 3982 3120 3991
rect 3144 3982 3153 3991
rect 3411 3982 3420 3991
rect 3444 3982 3453 3991
rect 3957 3982 3966 3991
rect 2157 3889 2166 3899
rect 3982 3980 3991 3989
rect 2511 3889 2520 3899
rect 3711 3964 3720 3973
rect 2157 3849 2166 3859
rect 2511 3849 2520 3859
rect 3982 3734 3991 3743
rect 1009 3711 1018 3720
rect 3982 3680 3991 3689
rect 3982 3647 3991 3656
rect 3850 3556 3860 3566
rect 3890 3556 3900 3566
rect 1009 3411 1018 3420
rect 1101 3411 1111 3420
rect 1141 3411 1151 3420
rect 3850 3380 3860 3389
rect 3890 3380 3900 3389
rect 3982 3380 3991 3389
rect 1009 3144 1018 3153
rect 1101 3144 1111 3153
rect 1141 3144 1151 3153
rect 1009 3057 1018 3066
rect 1101 3057 1111 3066
rect 1141 3057 1151 3066
rect 3850 2834 3860 2843
rect 3890 2834 3900 2843
rect 3982 2834 3991 2843
rect 1009 2811 1018 2820
rect 3982 2780 3991 2789
rect 3850 2534 3860 2543
rect 3890 2534 3900 2543
rect 3982 2534 3991 2543
rect 1009 2511 1018 2520
rect 1101 2511 1111 2520
rect 1141 2511 1151 2520
rect 3982 2480 3991 2489
rect 3850 2234 3860 2243
rect 3890 2234 3900 2243
rect 3982 2234 3991 2243
rect 1009 2211 1018 2220
rect 1101 2211 1111 2220
rect 1141 2211 1151 2220
rect 3982 2180 3991 2189
rect 3850 1934 3860 1943
rect 3890 1934 3900 1943
rect 3982 1934 3991 1943
rect 1009 1911 1018 1920
rect 1101 1911 1111 1920
rect 1141 1911 1151 1920
rect 3982 1880 3991 1889
rect 3850 1634 3860 1643
rect 3890 1634 3900 1643
rect 3982 1634 3991 1643
rect 1009 1611 1018 1620
rect 1101 1611 1111 1620
rect 1141 1611 1151 1620
rect 3982 1580 3991 1589
rect 3850 1334 3860 1343
rect 3890 1334 3900 1343
rect 3982 1334 3991 1343
rect 1009 1311 1018 1320
rect 1101 1311 1111 1320
rect 1141 1311 1151 1320
rect 3982 1280 3991 1289
rect 2645 1141 2655 1151
rect 1009 1044 1018 1053
rect 1311 1027 1320 1036
rect 1611 1027 1620 1036
rect 1911 1027 1920 1036
rect 2211 1027 2220 1036
rect 1026 1009 1035 1018
rect 1257 1009 1266 1018
rect 1557 1009 1566 1018
rect 1857 1009 1866 1018
rect 2157 1009 2166 1018
rect 2457 1009 2466 1018
rect 2811 1027 2820 1036
rect 3111 1027 3120 1036
rect 3411 1027 3420 1036
rect 3711 1027 3720 1036
rect 3982 1034 3991 1043
rect 3057 1009 3066 1018
rect 3357 1009 3366 1018
rect 3657 1009 3666 1018
rect 3957 1009 3966 1018
<< metal2 >>
rect 1020 4740 1274 4994
rect 1320 4740 1574 4994
rect 1620 4740 1874 4994
rect 1920 4740 2174 4994
rect 2220 4740 2474 4994
rect 2520 4740 2774 4994
rect 2820 4740 3074 4994
rect 3120 4740 3374 4994
rect 3420 4740 3674 4994
rect 3720 4740 3974 4994
rect 1011 3991 1020 4000
rect 1044 3991 1053 4000
rect 0 3720 254 3974
rect 1257 3973 1266 4000
rect 1311 3991 1320 4000
rect 1344 3991 1353 4000
rect 1557 3973 1566 4000
rect 1000 3957 1018 3966
rect 1257 3964 1309 3973
rect 1009 3955 1018 3957
rect 1009 3946 1301 3955
rect 1027 3928 1293 3937
rect 1000 3744 1018 3753
rect 1009 3720 1018 3744
rect 1000 3711 1009 3720
rect 0 3420 254 3674
rect 1027 3666 1036 3928
rect 1289 3879 1293 3928
rect 1297 3879 1301 3946
rect 1305 3879 1309 3964
rect 1400 3964 1566 3973
rect 1611 3973 1620 4000
rect 1400 3879 1404 3964
rect 1644 3955 1653 4000
rect 1857 3991 1866 4000
rect 1911 3973 1920 4000
rect 1453 3946 1653 3955
rect 1453 3879 1457 3946
rect 1944 3937 1953 4000
rect 2157 3991 2166 4000
rect 2511 3991 2520 4000
rect 2544 3991 2553 4000
rect 2520 3982 2544 3991
rect 1461 3928 1953 3937
rect 2757 3937 2766 4000
rect 2811 3991 2820 4000
rect 2844 3991 2853 4000
rect 3057 3955 3066 4000
rect 3111 3991 3120 4000
rect 3144 3991 3153 4000
rect 3357 3973 3366 4000
rect 3411 3991 3420 4000
rect 3444 3991 3453 4000
rect 3657 3991 3666 4000
rect 3503 3982 3666 3991
rect 3357 3964 3475 3973
rect 3057 3946 3467 3955
rect 2757 3928 3459 3937
rect 1461 3879 1465 3928
rect 2157 3859 2166 3889
rect 2511 3859 2520 3889
rect 3455 3879 3459 3928
rect 3463 3879 3467 3946
rect 3471 3879 3475 3964
rect 3503 3879 3507 3982
rect 3711 3973 3720 4000
rect 3744 3955 3753 4000
rect 3957 3991 3966 4000
rect 3991 3980 4000 3989
rect 3629 3946 3753 3955
rect 3982 3947 4000 3956
rect 3629 3879 3633 3946
rect 3982 3937 3991 3947
rect 3641 3928 3991 3937
rect 3641 3879 3645 3928
rect 3697 3906 3936 3915
rect 3697 3879 3701 3906
rect 3721 3888 3918 3897
rect 3721 3879 3725 3888
rect 1000 3657 1036 3666
rect 1065 3760 1121 3764
rect 1000 3444 1018 3453
rect 1009 3420 1018 3444
rect 1000 3411 1009 3420
rect 0 3120 254 3374
rect 1065 3366 1074 3760
rect 1000 3357 1074 3366
rect 1083 3750 1121 3754
rect 1000 3144 1009 3153
rect 1009 3120 1018 3144
rect 1000 3111 1018 3120
rect 0 2820 254 3074
rect 1000 3057 1009 3066
rect 1083 2853 1092 3750
rect 3860 3556 3890 3566
rect 1111 3411 1141 3420
rect 3860 3380 3890 3389
rect 1111 3144 1141 3153
rect 3909 3143 3918 3888
rect 3927 3443 3936 3906
rect 3991 3734 4000 3743
rect 4740 3720 4994 3974
rect 3991 3680 4000 3689
rect 3991 3647 4000 3656
rect 3927 3434 4000 3443
rect 4740 3420 4994 3674
rect 3991 3380 4000 3389
rect 3982 3356 3991 3380
rect 3982 3347 4000 3356
rect 3909 3134 4000 3143
rect 4740 3120 4994 3374
rect 3982 3080 4000 3089
rect 1111 3057 1141 3066
rect 1000 2844 1092 2853
rect 3982 3056 3991 3080
rect 3982 3047 4000 3056
rect 3982 2843 3991 3047
rect 3860 2834 3890 2843
rect 3991 2834 4000 2843
rect 4740 2820 4994 3074
rect 1000 2811 1009 2820
rect 3991 2780 4000 2789
rect 0 2520 254 2774
rect 1000 2757 1088 2766
rect 1000 2544 1018 2553
rect 1009 2520 1018 2544
rect 1000 2511 1009 2520
rect 0 2220 254 2474
rect 1000 2457 1075 2466
rect 1000 2244 1018 2253
rect 1009 2220 1018 2244
rect 1000 2211 1009 2220
rect 0 1920 254 2174
rect 1000 2157 1062 2166
rect 1000 1944 1018 1953
rect 1009 1920 1018 1944
rect 1000 1911 1009 1920
rect 0 1620 254 1874
rect 1000 1857 1049 1866
rect 1000 1644 1018 1653
rect 1009 1620 1018 1644
rect 1000 1611 1009 1620
rect 0 1320 254 1574
rect 1000 1557 1036 1566
rect 1027 1458 1036 1557
rect 1040 1473 1049 1857
rect 1053 1552 1062 2157
rect 1066 1560 1075 2457
rect 1079 1568 1088 2757
rect 3910 2747 4000 2756
rect 3860 2534 3890 2543
rect 1111 2511 1141 2520
rect 3860 2234 3890 2243
rect 1111 2211 1141 2220
rect 3860 1934 3890 1943
rect 1111 1911 1141 1920
rect 3910 1680 3919 2747
rect 3991 2534 4000 2543
rect 4740 2520 4994 2774
rect 3991 2480 4000 2489
rect 3880 1676 3919 1680
rect 3928 2447 4000 2456
rect 3860 1634 3890 1643
rect 1111 1611 1141 1620
rect 3928 1576 3937 2447
rect 3991 2234 4000 2243
rect 4740 2220 4994 2474
rect 3991 2180 4000 2189
rect 3880 1572 3937 1576
rect 3946 2147 4000 2156
rect 1079 1564 1121 1568
rect 3946 1563 3955 2147
rect 3991 1934 4000 1943
rect 4740 1920 4994 2174
rect 3991 1880 4000 1889
rect 1066 1556 1121 1560
rect 3880 1559 3955 1563
rect 3964 1847 4000 1856
rect 1053 1548 1121 1552
rect 3964 1550 3973 1847
rect 3991 1634 4000 1643
rect 4740 1620 4994 1874
rect 3991 1580 4000 1589
rect 3880 1546 3973 1550
rect 3982 1547 4000 1556
rect 1040 1469 1121 1473
rect 1416 1462 1420 1466
rect 3730 1462 3734 1466
rect 3982 1458 3991 1547
rect 1027 1454 1121 1458
rect 3880 1454 3991 1458
rect 1027 1446 1121 1450
rect 3880 1446 3973 1450
rect 1000 1344 1018 1353
rect 1009 1320 1018 1344
rect 1000 1311 1009 1320
rect 3 1023 257 1277
rect 1027 1266 1036 1446
rect 3860 1334 3890 1343
rect 1111 1311 1141 1320
rect 1000 1257 1036 1266
rect 3964 1256 3973 1446
rect 3991 1334 4000 1343
rect 4740 1320 4994 1574
rect 3991 1280 4000 1289
rect 3964 1247 4000 1256
rect 1300 1054 1308 1121
rect 1000 1044 1009 1053
rect 1009 1025 1018 1044
rect 1008 1024 1018 1025
rect 1044 1045 1308 1054
rect 1007 1023 1017 1024
rect 1006 1022 1016 1023
rect 1005 1021 1015 1022
rect 1004 1020 1014 1021
rect 1000 1019 1013 1020
rect 1000 1018 1012 1019
rect 1000 1017 1011 1018
rect 1024 1017 1026 1018
rect 1000 1016 1010 1017
rect 1023 1016 1026 1017
rect 1000 1015 1009 1016
rect 1022 1015 1026 1016
rect 1000 1014 1008 1015
rect 1021 1014 1026 1015
rect 1000 1013 1007 1014
rect 1020 1013 1026 1014
rect 1000 1012 1006 1013
rect 1019 1012 1026 1013
rect 1000 1011 1005 1012
rect 1018 1011 1026 1012
rect 1017 1010 1026 1011
rect 1016 1009 1026 1010
rect 1015 1008 1025 1009
rect 1014 1007 1024 1008
rect 1013 1006 1023 1007
rect 1012 1005 1022 1006
rect 1011 1004 1021 1005
rect 1011 1000 1020 1004
rect 1044 1000 1053 1045
rect 1257 1000 1266 1009
rect 1311 1000 1320 1027
rect 1454 1018 1462 1121
rect 1608 1054 1616 1121
rect 1762 1054 1770 1121
rect 1915 1072 1925 1121
rect 2645 1092 2655 1141
rect 2644 1091 2656 1092
rect 2643 1090 2657 1091
rect 2642 1089 2658 1090
rect 2641 1088 2659 1089
rect 2640 1087 2660 1088
rect 2639 1086 2661 1087
rect 2638 1085 2662 1086
rect 2637 1084 2663 1085
rect 2636 1083 2664 1084
rect 2635 1082 2665 1083
rect 2634 1081 2666 1082
rect 2633 1080 2667 1081
rect 2632 1079 2668 1080
rect 2631 1078 2669 1079
rect 2630 1077 2670 1078
rect 2629 1076 2671 1077
rect 2628 1075 2672 1076
rect 2627 1074 2673 1075
rect 2626 1073 2674 1074
rect 2625 1072 2675 1073
rect 1915 1063 2253 1072
rect 2624 1071 2676 1072
rect 2623 1070 2677 1071
rect 2622 1069 2678 1070
rect 2621 1068 2679 1069
rect 2620 1067 2680 1068
rect 2619 1066 2681 1067
rect 2618 1065 2682 1066
rect 3148 1065 3156 1121
rect 2617 1064 2683 1065
rect 2616 1063 2684 1064
rect 1608 1045 1653 1054
rect 1762 1045 1953 1054
rect 1344 1009 1462 1018
rect 1344 1000 1353 1009
rect 1557 1000 1566 1009
rect 1611 1000 1620 1027
rect 1644 1000 1653 1045
rect 1857 1000 1866 1009
rect 1911 1000 1920 1027
rect 1944 1000 1953 1045
rect 2157 1000 2166 1009
rect 2211 1000 2220 1027
rect 2244 1000 2253 1063
rect 2615 1062 2685 1063
rect 2614 1061 2686 1062
rect 2613 1060 2687 1061
rect 2612 1059 2688 1060
rect 2611 1058 2689 1059
rect 2610 1057 2690 1058
rect 2609 1056 2691 1057
rect 2844 1056 3156 1065
rect 2608 1055 2692 1056
rect 2607 1054 2693 1055
rect 2606 1053 2694 1054
rect 2605 1052 2695 1053
rect 2604 1051 2696 1052
rect 2603 1050 2697 1051
rect 2457 1000 2466 1009
rect 2602 1000 2698 1050
rect 2811 1000 2820 1027
rect 2844 1000 2853 1056
rect 3057 1000 3066 1009
rect 3111 1000 3120 1027
rect 3302 1018 3310 1121
rect 3144 1009 3310 1018
rect 3144 1000 3153 1009
rect 3357 1000 3366 1009
rect 3411 1000 3420 1027
rect 3456 1018 3464 1121
rect 3610 1076 3618 1121
rect 3610 1067 3753 1076
rect 3444 1009 3464 1018
rect 3444 1000 3453 1009
rect 3657 1000 3666 1009
rect 3711 1000 3720 1027
rect 3744 1000 3753 1067
rect 3991 1034 4000 1043
rect 4740 1020 4994 1274
rect 3957 1000 3966 1009
rect 1020 0 1274 254
rect 1320 0 1574 254
rect 1620 0 1874 254
rect 1920 0 2174 254
rect 2220 0 2474 254
rect 2520 0 2774 254
rect 2820 0 3074 254
rect 3120 0 3374 254
rect 3420 0 3674 254
rect 3720 0 3974 254
use logo  logo_0
timestamp 1383914834
transform 1 0 1490 0 1 3485
box 0 4 1940 292
use top  top_0
timestamp 1383913817
transform 1 0 1306 0 1 -905
box -185 2026 2574 4784
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1383894587
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< labels >>
rlabel metal2 1023 1257 1032 1266 0 D2
rlabel metal2 3720 0 3974 254 0 W15
rlabel metal2 3420 0 3674 254 0 W14
rlabel metal2 3120 0 3374 254 0 W13
rlabel metal2 2820 0 3074 254 0 W12
rlabel metal2 2520 0 2774 254 0 GND
rlabel metal2 2220 0 2474 254 0 W4
rlabel metal2 1920 0 2174 254 0 W3
rlabel metal2 1620 0 1874 254 0 W2
rlabel metal2 1320 0 1574 254 0 W1
rlabel metal2 1020 0 1274 254 0 W0
rlabel metal2 4740 3720 4994 3974 0 TFQ
rlabel metal2 4740 3420 4994 3674 0 TFD
rlabel metal2 4740 3120 4994 3374 0 TFC
rlabel metal2 4740 2820 4994 3074 0 NC
rlabel metal2 4740 2520 4994 2774 0 PCLKO
rlabel metal2 4740 2220 4994 2474 0 PSO
rlabel metal2 4740 1920 4994 2174 0 TESTO
rlabel metal2 4740 1620 4994 1874 0 SO
rlabel metal2 4740 1320 4994 1574 0 LDO
rlabel metal2 4740 1020 4994 1274 0 SCLKO
rlabel metal2 1020 4740 1274 4994 0 TPZI
rlabel metal2 1320 4740 1574 4994 0 TPWI
rlabel metal2 1620 4740 1874 4994 0 TPZO
rlabel metal2 1920 4740 2174 4994 0 TPQO
rlabel metal2 2220 4740 2474 4994 0 VDD
rlabel metal2 2520 4740 2774 4994 0 TSSI
rlabel metal2 2820 4740 3074 4994 0 TSLDI
rlabel metal2 3120 4740 3374 4994 0 TSCI
rlabel metal2 3420 4740 3674 4994 0 TSZ
rlabel metal2 3720 4740 3974 4994 0 TSSO
rlabel metal2 0 1320 254 1574 0 LDI
rlabel metal2 0 1620 254 1874 0 SI
rlabel metal2 0 1920 254 2174 0 TESTI
rlabel metal2 0 2220 254 2474 0 PSI
rlabel metal2 0 2520 254 2774 0 PCLKI
rlabel metal2 0 2820 254 3074 0 TIO
rlabel metal2 0 3120 254 3374 0 TII
rlabel metal2 0 3420 254 3674 0 TPQI
rlabel metal2 0 3720 254 3974 0 TPCI
rlabel metal2 3 1023 257 1277 0 SCLKI
rlabel metal2 3730 1462 3734 1466 0 D_SSO
rlabel metal2 3882 1446 3892 1450 0 D_SCLKO
rlabel metal2 1104 1469 1111 1473 0 D_SI
rlabel metal2 1416 1462 1420 1466 0 D_SQ0
<< end >>
