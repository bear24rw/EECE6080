magic
tech scmos
timestamp 1380590399
<< ntransistor >>
rect -53 33 -51 37
rect -37 33 -35 37
rect -21 33 -19 37
rect -5 33 -3 37
rect 11 33 13 37
rect 27 33 29 37
rect -45 13 -43 17
rect -13 13 -11 17
rect 43 33 45 37
rect 35 13 37 17
rect -53 -45 -51 -41
rect -37 -45 -35 -41
rect -21 -45 -19 -41
rect -5 -45 -3 -41
rect 11 -45 13 -41
rect 27 -45 29 -41
rect 43 -45 45 -41
<< ptransistor >>
rect -53 49 -51 53
rect -37 49 -35 53
rect -21 49 -19 53
rect -5 49 -3 53
rect 11 49 13 53
rect 27 49 29 53
rect 43 49 45 53
rect -45 -3 -43 1
rect -13 -3 -11 1
rect 35 -3 37 1
rect -53 -29 -51 -25
rect -37 -29 -35 -25
rect -21 -29 -19 -25
rect -5 -29 -3 -25
rect 11 -29 13 -25
rect 27 -29 29 -25
rect 43 -29 45 -25
<< ndiffusion >>
rect -54 33 -53 37
rect -51 33 -50 37
rect -38 33 -37 37
rect -35 33 -34 37
rect -22 33 -21 37
rect -19 33 -18 37
rect -6 33 -5 37
rect -3 33 -2 37
rect 10 33 11 37
rect 13 33 14 37
rect 26 33 27 37
rect 29 33 30 37
rect -46 13 -45 17
rect -43 13 -42 17
rect -14 13 -13 17
rect -11 13 -10 17
rect 42 33 43 37
rect 45 33 46 37
rect 34 13 35 17
rect 37 13 38 17
rect -54 -45 -53 -41
rect -51 -45 -37 -41
rect -35 -45 -34 -41
rect -22 -45 -21 -41
rect -19 -45 -18 -41
rect -6 -45 -5 -41
rect -3 -45 11 -41
rect 13 -45 14 -41
rect 26 -45 27 -41
rect 29 -45 43 -41
rect 45 -45 46 -41
<< pdiffusion >>
rect -54 49 -53 53
rect -51 49 -50 53
rect -38 49 -37 53
rect -35 49 -34 53
rect -22 49 -21 53
rect -19 49 -18 53
rect -6 49 -5 53
rect -3 49 -2 53
rect 10 49 11 53
rect 13 49 14 53
rect 26 49 27 53
rect 29 49 30 53
rect 42 49 43 53
rect 45 49 46 53
rect -46 -3 -45 1
rect -43 -3 -42 1
rect -14 -3 -13 1
rect -11 -3 -10 1
rect 34 -3 35 1
rect 37 -3 38 1
rect -54 -29 -53 -25
rect -51 -29 -50 -25
rect -38 -29 -37 -25
rect -35 -29 -34 -25
rect -22 -29 -21 -25
rect -19 -29 -18 -25
rect -6 -29 -5 -25
rect -3 -29 -2 -25
rect 10 -29 11 -25
rect 13 -29 14 -25
rect 26 -29 27 -25
rect 29 -29 30 -25
rect 42 -29 43 -25
rect 45 -29 46 -25
<< ndcontact >>
rect -58 33 -54 37
rect -50 33 -46 37
rect -42 33 -38 37
rect -34 33 -30 37
rect -26 33 -22 37
rect -18 33 -14 37
rect -10 33 -6 37
rect -2 33 2 37
rect 6 33 10 37
rect 14 33 18 37
rect 22 33 26 37
rect 30 33 34 37
rect -50 13 -46 17
rect -42 13 -38 17
rect -18 13 -14 17
rect -10 13 -6 17
rect 38 33 42 37
rect 46 33 50 37
rect 30 13 34 17
rect 38 13 42 17
rect -58 -45 -54 -41
rect -34 -45 -30 -41
rect -26 -45 -22 -41
rect -18 -45 -14 -41
rect -10 -45 -6 -41
rect 14 -45 18 -41
rect 22 -45 26 -41
rect 46 -45 50 -41
<< pdcontact >>
rect -58 49 -54 53
rect -50 49 -46 53
rect -42 49 -38 53
rect -34 49 -30 53
rect -26 49 -22 53
rect -18 49 -14 53
rect -10 49 -6 53
rect -2 49 2 53
rect 6 49 10 53
rect 14 49 18 53
rect 22 49 26 53
rect 30 49 34 53
rect 38 49 42 53
rect 46 49 50 53
rect -50 -3 -46 1
rect -42 -3 -38 1
rect -18 -3 -14 1
rect -10 -3 -6 1
rect 30 -3 34 1
rect 38 -3 42 1
rect -58 -29 -54 -25
rect -50 -29 -46 -25
rect -42 -29 -38 -25
rect -34 -29 -30 -25
rect -26 -29 -22 -25
rect -18 -29 -14 -25
rect -10 -29 -6 -25
rect -2 -29 2 -25
rect 6 -29 10 -25
rect 14 -29 18 -25
rect 22 -29 26 -25
rect 30 -29 34 -25
rect 38 -29 42 -25
rect 46 -29 50 -25
<< polysilicon >>
rect -53 66 -51 70
rect -53 53 -51 62
rect -37 53 -35 55
rect -21 53 -19 55
rect -5 53 -3 55
rect 11 53 13 70
rect 27 53 29 55
rect 43 53 45 62
rect -53 37 -51 49
rect -53 -25 -51 33
rect -45 17 -43 41
rect -37 37 -35 49
rect -21 37 -19 49
rect -5 45 -3 49
rect -37 24 -35 33
rect -21 24 -19 33
rect -13 17 -11 41
rect -5 37 -3 41
rect 11 37 13 49
rect 27 45 29 49
rect 27 37 29 41
rect -5 31 -3 33
rect -45 1 -43 13
rect -13 1 -11 13
rect -45 -5 -43 -3
rect -13 -5 -11 -3
rect -37 -25 -35 -23
rect -21 -25 -19 -16
rect -5 -25 -3 -16
rect 11 -25 13 33
rect 27 31 29 33
rect 35 17 37 41
rect 43 37 45 49
rect 43 31 45 33
rect 35 1 37 13
rect 35 -5 37 -3
rect 27 -25 29 -23
rect 43 -25 45 -23
rect -53 -41 -51 -29
rect -37 -33 -35 -29
rect -37 -41 -35 -37
rect -21 -41 -19 -29
rect -5 -41 -3 -29
rect 11 -41 13 -29
rect 27 -33 29 -29
rect 27 -41 29 -37
rect 43 -41 45 -29
rect -53 -47 -51 -45
rect -37 -47 -35 -45
rect -21 -47 -19 -45
rect -5 -47 -3 -45
rect 11 -47 13 -45
rect 27 -47 29 -45
rect 43 -54 45 -45
<< polycontact >>
rect -54 62 -50 66
rect 42 62 46 66
rect -46 41 -42 45
rect -14 41 -10 45
rect -6 41 -2 45
rect -38 20 -34 24
rect -22 20 -18 24
rect 26 41 30 45
rect 34 41 38 45
rect -22 -16 -18 -12
rect -6 -16 -2 -12
rect -38 -37 -34 -33
rect 26 -37 30 -33
rect 42 -58 46 -54
<< metal1 >>
rect -50 62 42 66
rect -62 56 58 59
rect -58 53 -54 56
rect -34 53 -30 56
rect -46 45 -42 53
rect -26 53 -22 56
rect -2 53 2 56
rect 14 53 18 56
rect -14 45 -10 53
rect 22 53 26 56
rect 46 53 50 56
rect 6 45 10 49
rect 34 45 38 53
rect -58 41 -46 45
rect -26 41 -14 45
rect -2 41 26 45
rect 38 41 50 45
rect -58 37 -54 41
rect -26 37 -22 41
rect 6 37 10 41
rect 46 37 50 41
rect -46 33 -42 37
rect -14 33 -10 37
rect 34 33 38 37
rect -34 30 -30 33
rect -2 30 2 33
rect 22 30 26 33
rect -62 27 58 30
rect -58 20 -38 24
rect -34 20 -22 24
rect -58 9 -54 20
rect 38 17 42 27
rect -62 5 -54 9
rect -38 13 -18 17
rect -6 13 30 17
rect -50 9 -46 13
rect -50 5 58 9
rect -50 1 -46 5
rect -18 1 -14 5
rect 30 1 34 5
rect -42 -6 -38 -3
rect -10 -6 -6 -3
rect 38 -6 42 -3
rect -62 -9 58 -6
rect -62 -16 -22 -12
rect -18 -16 -6 -12
rect -2 -16 58 -12
rect -62 -22 58 -19
rect -58 -25 -54 -22
rect -34 -25 -30 -22
rect -18 -25 -14 -22
rect 14 -25 18 -22
rect -46 -33 -42 -25
rect -26 -33 -22 -29
rect 2 -33 6 -25
rect 22 -25 26 -22
rect 46 -25 50 -22
rect 34 -33 38 -25
rect -58 -37 -42 -33
rect -34 -37 -22 -33
rect -58 -41 -54 -37
rect -26 -41 -22 -37
rect -10 -37 26 -33
rect 34 -37 59 -33
rect -10 -41 -6 -37
rect 46 -41 50 -37
rect -58 -54 -54 -45
rect -34 -48 -30 -45
rect -18 -48 -14 -45
rect 14 -48 18 -45
rect 22 -48 26 -45
rect -34 -51 52 -48
rect -58 -58 42 -54
rect 49 -61 52 -51
rect 55 -58 59 -37
rect -61 -65 59 -61
<< labels >>
rlabel metal1 -62 56 -58 59 0 VDD
rlabel metal1 -62 27 -58 30 0 GND
rlabel metal1 -62 5 -58 9 0 C_IN
rlabel metal1 -62 -9 -58 -6 0 VDD
rlabel metal1 -62 -16 -58 -12 0 S
rlabel metal1 -62 -22 -58 -19 0 VDD
rlabel metal1 -61 -65 -58 -61 0 GND
rlabel metal1 55 -58 59 -54 0 F
rlabel metal1 50 5 58 9 0 C_OUT
rlabel polysilicon -53 66 -51 70 0 B
rlabel polysilicon 11 66 13 70 0 A
<< end >>
