magic
tech scmos
timestamp 1383821139
<< metal1 >>
rect -17 109 2446 113
rect 2442 80 2446 109
rect -13 36 -9 40
<< m2contact >>
rect 10 117 14 121
rect -21 109 -17 113
rect 2438 80 2442 84
rect 10 1 14 5
<< metal2 >>
rect -21 196 6 200
rect -21 113 -17 196
rect 10 121 14 128
rect 101 93 105 129
rect 253 93 257 129
rect 405 93 409 129
rect 557 93 561 129
rect 709 93 713 129
rect 861 93 865 129
rect 1013 93 1017 129
rect 1165 93 1169 129
rect 1317 93 1321 129
rect 1469 93 1473 129
rect 1621 93 1625 129
rect 1773 93 1777 129
rect 1925 93 1929 129
rect 2077 93 2081 129
rect 2229 93 2233 129
rect 2381 93 2385 129
rect 10 5 14 16
<< end >>
