magic
tech scmos
timestamp 1381994511
use MUX2X1  MUX2X1_0
timestamp 1053021328
transform 1 0 5 0 1 3
box -5 -3 53 105
use DFFPOSX1  DFFPOSX1_0
timestamp 1048618183
transform 1 0 47 0 1 3
box -8 -3 104 105
<< end >>
