magic
tech scmos
timestamp 1383875311
<< nwell >>
rect -7 48 39 105
<< ntransistor >>
rect 10 6 12 26
rect 15 6 17 26
rect 23 6 25 16
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 9 6 10 26
rect 12 6 15 26
rect 17 6 18 26
rect 22 6 23 16
rect 25 6 26 16
<< pdiffusion >>
rect 6 57 7 94
rect 2 54 7 57
rect 9 60 10 94
rect 14 60 15 94
rect 9 54 15 60
rect 17 54 18 94
rect 22 54 23 94
rect 25 54 26 94
<< ndcontact >>
rect 5 6 9 26
rect 18 6 22 26
rect 26 6 30 16
<< pdcontact >>
rect 2 57 6 94
rect 10 60 14 94
rect 18 54 22 94
rect 26 54 30 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect 0 98 4 102
rect 18 98 22 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 49 9 54
rect 4 29 6 47
rect 15 41 17 54
rect 14 37 17 41
rect 4 27 12 29
rect 10 26 12 27
rect 15 26 17 37
rect 23 16 25 54
rect 10 4 12 6
rect 15 4 17 6
rect 23 4 25 6
<< polycontact >>
rect 6 45 10 49
rect 10 37 14 41
rect 25 19 29 23
<< metal1 >>
rect -2 102 34 103
rect -2 98 0 102
rect 4 98 18 102
rect 22 98 34 102
rect -2 97 34 98
rect 10 94 14 97
rect 2 54 18 57
rect 2 45 6 47
rect 26 47 29 54
rect 2 44 10 45
rect 18 44 30 47
rect 2 43 6 44
rect 10 33 14 37
rect 18 26 21 44
rect 26 23 30 27
rect 5 3 9 6
rect 26 3 30 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< m1p >>
rect 2 43 6 47
rect 26 43 30 47
rect 10 33 14 37
rect 26 23 30 27
<< labels >>
rlabel metal1 4 0 4 0 1 gnd
rlabel metal1 4 100 4 100 5 vdd
rlabel metal1 4 45 4 45 1 A
rlabel metal1 12 35 12 35 1 B
rlabel metal1 28 45 28 45 1 Y
rlabel metal1 28 25 28 25 1 C
<< end >>
