magic
tech scmos
timestamp 1380848338
<< polysilicon >>
rect 8 135 10 139
rect 72 135 74 139
rect 128 135 130 139
rect 192 135 194 139
rect 248 135 250 139
rect 312 135 314 139
<< metal1 >>
rect -3 70 0 74
rect 360 70 367 74
rect 363 53 367 70
rect 360 49 367 53
rect 116 11 120 15
rect 236 11 240 15
rect 356 11 360 15
use slice  slice_0
array 0 2 120 0 0 135
timestamp 1380769700
transform 1 0 61 0 1 65
box -61 -65 59 70
<< labels >>
rlabel polysilicon 8 135 10 139 0 B0
rlabel polysilicon 72 135 74 139 0 A0
rlabel polysilicon 128 135 130 139 0 B1
rlabel polysilicon 192 135 194 139 0 A1
rlabel polysilicon 248 135 250 139 0 B2
rlabel polysilicon 312 135 314 139 0 A2
rlabel metal1 -3 70 0 74 0 GND
rlabel metal1 116 11 120 15 0 F0
rlabel metal1 236 11 240 15 0 F1
rlabel metal1 356 11 360 15 0 F2
<< end >>
