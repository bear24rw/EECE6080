magic
tech scmos
timestamp 1383010634
<< metal2 >>
rect 22 -83 26 4
rect 183 -77 187 4
rect 344 -71 348 4
rect 505 -65 509 4
rect 666 -59 670 4
rect 827 -53 831 4
rect 988 -47 992 4
rect 1149 -41 1153 4
rect 1310 -35 1314 4
rect 1471 -29 1475 4
rect 1632 -23 1636 4
rect 1793 -17 1797 4
rect 1954 -11 1958 4
rect 2115 -5 2119 4
rect 2276 1 2280 4
rect 2276 -2 2405 1
rect 2115 -8 2405 -5
rect 1954 -14 2405 -11
rect 1793 -20 2405 -17
rect 1631 -26 2405 -23
rect 1471 -32 2405 -29
rect 1310 -38 2405 -35
rect 1149 -44 2405 -41
rect 988 -50 2405 -47
rect 827 -56 2405 -53
rect 666 -62 2405 -59
rect 505 -68 2405 -65
rect 344 -74 2405 -71
rect 183 -80 2405 -77
rect 22 -86 2405 -83
use shift_slice  shift_slice_0
array 0 14 161 0 0 107
timestamp 1382932048
transform 1 0 0 0 1 4
box -17 0 151 108
<< end >>
