magic
tech scmos
timestamp 1382939220
<< metal1 >>
rect -1 162 3 165
rect -8 153 -1 156
rect -1 109 2289 113
rect 2293 109 2343 113
rect 2 0 6 12
<< m2contact >>
rect -5 161 -1 165
rect -12 152 -8 156
rect -5 109 -1 113
rect 2343 109 2347 113
rect 2 12 6 16
<< metal2 >>
rect -12 40 -8 152
rect -5 113 -1 161
rect 101 93 105 129
rect 257 93 261 129
rect 413 93 417 129
rect 569 93 573 129
rect 725 93 729 129
rect 881 93 885 129
rect 1037 93 1041 129
rect 1193 93 1197 129
rect 1349 93 1353 129
rect 1505 93 1509 129
rect 1661 93 1665 129
rect 1817 93 1821 129
rect 1973 93 1977 129
rect 2129 93 2133 129
rect 2285 93 2289 129
rect 2343 49 2347 109
<< end >>
