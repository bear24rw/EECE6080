magic
tech scmos
timestamp 1383894587
<< polysilicon >>
rect 0 0 150 2900
<< end >>
