magic
tech scmos
timestamp 1383882935
<< metal2 >>
rect 2018 1819 2121 1823
rect -449 5 -445 1785
rect 2018 1751 2114 1755
rect 2018 1635 2108 1639
rect 2018 1519 2102 1523
rect 2018 1403 2096 1407
rect 2018 1287 2090 1291
rect 2018 1171 2084 1175
rect 2018 1055 2078 1059
rect 2018 939 2072 943
rect 2018 823 2066 827
rect 2018 707 2060 711
rect 2018 591 2054 595
rect 2018 475 2048 479
rect 2018 359 2042 363
rect 2018 243 2036 247
rect 2018 127 2030 131
rect -440 79 -414 83
rect -440 5 -436 79
rect 2027 -1 2030 127
rect 2033 -1 2036 243
rect 2039 -1 2042 359
rect 2045 -1 2048 475
rect 2051 -1 2054 591
rect 2057 -1 2060 707
rect 2063 -1 2066 823
rect 2069 -1 2072 939
rect 2075 -1 2078 1055
rect 2081 -1 2084 1171
rect 2087 -1 2090 1287
rect 2093 -1 2096 1403
rect 2099 -1 2102 1519
rect 2105 -1 2108 1635
rect 2111 -1 2114 1751
rect 2117 -1 2121 1819
use pin_row_connect  pin_row_connect_0
array 0 0 2427 0 14 116
timestamp 1383821139
transform 1 0 -420 0 1 -1
box -21 1 2446 200
use pin_buffer  pin_buffer_0
array 0 0 46 0 15 116
timestamp 1383808422
transform 1 0 -460 0 1 -1
box 0 0 46 108
use pin_slice  pin_slice_0
array 0 15 152 0 15 116
timestamp 1383875311
transform 1 0 -324 0 1 112
box -100 -113 68 -5
use pin_testmode_mux  pin_testmode_mux_0
timestamp 1383816218
transform 1 0 -456 0 -1 5
box 0 0 131 108
<< end >>
