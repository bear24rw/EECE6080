magic
tech scmos
timestamp 1383821139
use top  top_0
timestamp 1383821139
transform 1 0 1315 0 1 -696
box -155 2193 2568 4477
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1072203966
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< end >>
