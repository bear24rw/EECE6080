magic
tech scmos
timestamp 1383634647
<< m2contact >>
rect 2402 50 2406 54
rect 2410 50 2414 54
<< metal2 >>
rect 2402 94 2406 110
rect 2409 87 2413 110
rect 2405 83 2413 87
rect 2416 61 2420 110
rect 2405 57 2420 61
rect 2410 54 2414 57
rect 2402 47 2406 50
rect 2423 47 2427 110
rect 2402 43 2427 47
rect 22 -83 26 4
rect 183 -77 187 4
rect 344 -71 348 4
rect 505 -65 509 4
rect 666 -59 670 4
rect 827 -53 831 4
rect 988 -47 992 4
rect 1149 -41 1153 4
rect 1310 -35 1314 4
rect 1471 -29 1475 4
rect 1632 -23 1636 4
rect 1793 -17 1797 4
rect 1954 -11 1958 4
rect 2115 -5 2119 4
rect 2276 1 2280 4
rect 2276 -2 2440 1
rect 2115 -8 2440 -5
rect 1954 -14 2440 -11
rect 1793 -20 2440 -17
rect 1631 -26 2440 -23
rect 1471 -32 2440 -29
rect 1310 -38 2440 -35
rect 1149 -44 2440 -41
rect 988 -50 2440 -47
rect 827 -56 2440 -53
rect 666 -62 2440 -59
rect 505 -68 2440 -65
rect 344 -74 2440 -71
rect 183 -80 2440 -77
rect 22 -86 2440 -83
use shift_slice  shift_slice_0
array 0 14 161 0 0 107
timestamp 1383629942
transform 1 0 0 0 1 4
box -17 0 151 108
use MUX2X1  MUX2X1_0
timestamp 1383629942
transform 1 0 2400 0 1 7
box -5 -3 53 105
<< end >>
