magic
tech scmos
timestamp 1383649547
<< error_s >>
rect 1195 1895 1199 1899
rect 1199 1869 1200 1887
rect 1217 1871 1219 1894
rect 1220 1891 1222 1893
rect 1220 1890 1224 1891
rect 1220 1871 1227 1890
rect 1198 1866 1200 1869
rect 1201 1840 1203 1866
rect 1220 1853 1224 1871
rect 1220 1845 1222 1853
rect 1201 1818 1203 1836
rect 1223 1833 1225 1840
rect 1220 1825 1222 1831
rect 1220 1820 1224 1825
rect 1199 1807 1200 1817
rect 1215 1816 1224 1820
rect 1220 1812 1224 1816
rect 1217 1805 1219 1812
rect 1220 1807 1227 1812
rect 1223 1803 1227 1807
rect 1195 1795 1199 1799
rect 1198 1765 1200 1769
rect 1198 1702 1200 1714
rect 1202 1706 1204 1710
rect 1198 1665 1200 1669
use INVX1  INVX1_0
timestamp 1383629942
transform 1 0 1213 0 1 1797
box -9 -3 26 105
use top  top_0
timestamp 1383649547
transform 1 0 1364 0 1 1679
box -198 -129 2445 1869
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1072203966
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< end >>
