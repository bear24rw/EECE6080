magic
tech scmos
timestamp 1383010634
<< metal2 >>
rect 2347 1636 2435 1640
rect 2347 1520 2429 1524
rect 2347 1404 2423 1408
rect 2347 1288 2417 1292
rect 2347 1172 2411 1176
rect 2347 1056 2405 1060
rect 2347 940 2399 944
rect 2347 824 2393 828
rect 2347 708 2387 712
rect 2347 592 2381 596
rect 2347 476 2375 480
rect 2347 360 2369 364
rect 2347 244 2363 248
rect 2347 128 2357 132
rect 2347 12 2351 16
rect 2348 0 2351 12
rect 2354 0 2357 128
rect 2360 0 2363 244
rect 2366 0 2369 360
rect 2372 0 2375 476
rect 2378 0 2381 592
rect 2384 0 2387 708
rect 2390 0 2393 824
rect 2396 0 2399 940
rect 2402 0 2405 1056
rect 2408 0 2411 1172
rect 2414 0 2417 1288
rect 2420 0 2423 1404
rect 2426 0 2429 1520
rect 2432 0 2435 1636
use pin_row_connect  pin_row_connect_0
array 0 0 98 0 13 116
timestamp 1382939220
transform 1 0 4 0 1 0
box -12 0 2347 165
use pin_slice  pin_slice_0
array 0 14 156 0 14 116
timestamp 1383010634
transform 1 0 100 0 1 113
box -100 -113 68 -5
<< end >>
