magic
tech scmos
timestamp 1383822934
<< nwell >>
rect -9 56 3 57
<< metal1 >>
rect -16 100 151 106
rect 45 45 60 49
rect 64 45 85 46
rect -16 0 151 6
<< m2contact >>
rect -9 46 -5 50
rect -1 46 3 50
rect 23 46 27 50
rect 137 46 141 50
rect 57 36 61 40
<< metal2 >>
rect 6 80 124 84
rect -9 53 3 57
rect -1 50 3 53
rect -9 42 -5 46
rect 6 42 10 80
rect -9 38 10 42
rect 15 54 35 58
rect 15 34 19 54
rect -9 30 19 34
rect 23 0 27 46
rect 31 16 35 54
rect 120 42 124 80
rect 137 57 141 106
rect 137 53 145 57
rect 137 50 141 53
rect 120 38 145 42
rect 57 16 61 36
rect 120 30 145 34
rect 120 16 124 30
rect 31 12 124 16
use mux  mux_0
timestamp 1383808422
transform 1 0 -16 0 1 0
box 0 0 73 108
use DFFPOSX1  DFFPOSX1_0
timestamp 1383803179
transform 1 0 47 0 1 3
box -8 -3 104 105
<< labels >>
rlabel metal1 145 100 151 106 0 VDD
rlabel metal1 145 0 151 6 0 GND
rlabel metal2 141 53 145 57 0 SO
rlabel metal2 23 0 27 6 0 Z
rlabel metal2 -9 38 -5 42 0 LDI
rlabel metal2 -9 30 -5 34 0 SCLKI
rlabel metal2 -9 53 -4 57 0 SI
<< end >>
