magic
tech scmos
timestamp 1383823585
<< nwell >>
rect 2366 2472 2378 2476
rect 2428 2464 2431 2468
rect 2434 2457 2436 2474
rect 2428 2451 2431 2455
rect 2434 2453 2436 2456
<< metal1 >>
rect -155 4469 2568 4477
rect -155 4367 -147 4469
rect -155 4361 -154 4367
rect -148 4361 -147 4367
rect -155 4251 -147 4361
rect -155 4245 -154 4251
rect -148 4245 -147 4251
rect -155 4135 -147 4245
rect -155 4129 -154 4135
rect -148 4129 -147 4135
rect -155 4019 -147 4129
rect -155 4013 -154 4019
rect -148 4013 -147 4019
rect -155 3903 -147 4013
rect -155 3897 -154 3903
rect -148 3897 -147 3903
rect -155 3787 -147 3897
rect -155 3781 -154 3787
rect -148 3781 -147 3787
rect -155 3671 -147 3781
rect -155 3665 -154 3671
rect -148 3665 -147 3671
rect -155 3555 -147 3665
rect -155 3549 -154 3555
rect -148 3549 -147 3555
rect -155 3439 -147 3549
rect -155 3433 -154 3439
rect -148 3433 -147 3439
rect -155 3323 -147 3433
rect -155 3317 -154 3323
rect -148 3317 -147 3323
rect -155 3207 -147 3317
rect -155 3201 -154 3207
rect -148 3201 -147 3207
rect -155 3091 -147 3201
rect -155 3085 -154 3091
rect -148 3085 -147 3091
rect -155 2975 -147 3085
rect -155 2969 -154 2975
rect -148 2969 -147 2975
rect -155 2859 -147 2969
rect -155 2853 -154 2859
rect -148 2853 -147 2859
rect -155 2743 -147 2853
rect -155 2737 -154 2743
rect -148 2737 -147 2743
rect -155 2627 -147 2737
rect -155 2621 -154 2627
rect -148 2621 -147 2627
rect -155 2427 -147 2621
rect -155 2421 -154 2427
rect -148 2421 -147 2427
rect -155 2201 -147 2421
rect -139 4453 2552 4461
rect -139 2217 -131 4453
rect -119 4361 -40 4367
rect 2544 4267 2552 4453
rect 2431 4261 2552 4267
rect -119 4245 -40 4251
rect 2544 4151 2552 4261
rect 2431 4145 2552 4151
rect -119 4129 -40 4135
rect 2544 4035 2552 4145
rect 2431 4029 2552 4035
rect -119 4013 -40 4019
rect 2544 3919 2552 4029
rect 2431 3913 2552 3919
rect -119 3897 -40 3903
rect 2544 3803 2552 3913
rect 2431 3797 2552 3803
rect -119 3781 -40 3787
rect 2544 3687 2552 3797
rect 2431 3681 2552 3687
rect -119 3665 -40 3671
rect 2544 3571 2552 3681
rect 2431 3565 2552 3571
rect -119 3549 -40 3555
rect 2544 3455 2552 3565
rect 2431 3449 2552 3455
rect -119 3433 -40 3439
rect 2544 3339 2552 3449
rect 2431 3333 2552 3339
rect -119 3317 -40 3323
rect 2544 3223 2552 3333
rect 2431 3217 2552 3223
rect -119 3201 -40 3207
rect 2544 3107 2552 3217
rect 2431 3101 2552 3107
rect -119 3085 -40 3091
rect 2544 2991 2552 3101
rect 2431 2985 2552 2991
rect -119 2969 -40 2975
rect 2544 2875 2552 2985
rect 2431 2869 2552 2875
rect -119 2853 -40 2859
rect 2544 2759 2552 2869
rect 2431 2753 2552 2759
rect -119 2737 -40 2743
rect 2544 2643 2552 2753
rect 2431 2637 2552 2643
rect -119 2621 -40 2627
rect 2432 2581 2537 2585
rect 2544 2527 2552 2637
rect 2431 2521 2552 2527
rect 2420 2487 2541 2491
rect 83 2480 2346 2484
rect 2358 2480 2374 2484
rect 2431 2477 2530 2481
rect 83 2472 2362 2476
rect 83 2464 2354 2468
rect 2362 2442 2366 2472
rect 2431 2464 2530 2468
rect 2537 2455 2541 2487
rect 2431 2451 2530 2455
rect -119 2421 -40 2427
rect 2431 2359 2537 2363
rect 2431 2351 2537 2355
rect 2544 2327 2552 2521
rect 2434 2321 2552 2327
rect 2544 2217 2552 2321
rect -139 2209 2552 2217
rect 2560 2201 2568 4469
rect -155 2193 2568 2201
<< m2contact >>
rect -154 4361 -148 4367
rect -154 4245 -148 4251
rect -154 4129 -148 4135
rect -154 4013 -148 4019
rect -154 3897 -148 3903
rect -154 3781 -148 3787
rect -154 3665 -148 3671
rect -154 3549 -148 3555
rect -154 3433 -148 3439
rect -154 3317 -148 3323
rect -154 3201 -148 3207
rect -154 3085 -148 3091
rect -154 2969 -148 2975
rect -154 2853 -148 2859
rect -154 2737 -148 2743
rect -154 2621 -148 2627
rect -154 2421 -148 2427
rect -125 4361 -119 4367
rect -125 4245 -119 4251
rect -125 4129 -119 4135
rect -125 4013 -119 4019
rect -125 3897 -119 3903
rect -125 3781 -119 3787
rect -125 3665 -119 3671
rect -125 3549 -119 3555
rect -125 3433 -119 3439
rect -125 3317 -119 3323
rect -125 3201 -119 3207
rect -125 3085 -119 3091
rect -125 2969 -119 2975
rect -125 2853 -119 2859
rect -125 2737 -119 2743
rect -125 2621 -119 2627
rect 2428 2581 2432 2585
rect 2537 2581 2541 2585
rect 79 2480 83 2484
rect 2346 2480 2350 2484
rect 2354 2480 2358 2484
rect 2378 2477 2382 2481
rect 2402 2477 2406 2481
rect 2427 2477 2431 2481
rect 2530 2477 2534 2481
rect 79 2472 83 2476
rect 2362 2472 2366 2476
rect 79 2464 83 2468
rect 2354 2464 2358 2468
rect 2427 2464 2431 2468
rect 2530 2464 2534 2468
rect 2427 2451 2431 2455
rect 2530 2451 2534 2455
rect 2537 2451 2541 2455
rect 2362 2438 2366 2442
rect -125 2421 -119 2427
rect 2427 2359 2431 2363
rect 2537 2359 2541 2363
rect 2427 2351 2431 2355
rect 2537 2351 2541 2355
<< metal2 >>
rect -148 4361 -125 4367
rect -148 4245 -125 4251
rect -148 4129 -125 4135
rect -148 4013 -125 4019
rect -148 3897 -125 3903
rect -148 3781 -125 3787
rect -148 3665 -125 3671
rect -148 3549 -125 3555
rect -148 3433 -125 3439
rect -148 3317 -125 3323
rect -148 3201 -125 3207
rect -148 3085 -125 3091
rect -148 2969 -125 2975
rect -148 2853 -125 2859
rect -148 2737 -125 2743
rect -148 2621 -125 2627
rect 2541 2581 2568 2585
rect 2431 2533 2437 2537
rect 76 2480 79 2484
rect 94 2476 98 2530
rect 246 2476 250 2530
rect 398 2476 402 2530
rect 550 2476 554 2530
rect 702 2476 706 2530
rect 854 2476 858 2530
rect 1006 2476 1010 2530
rect 1158 2476 1162 2530
rect 1310 2476 1314 2530
rect 1462 2476 1466 2530
rect 1614 2476 1618 2530
rect 1766 2476 1770 2530
rect 1918 2476 1922 2530
rect 2070 2476 2074 2530
rect 2222 2476 2226 2530
rect 2374 2492 2378 2530
rect 2374 2488 2382 2492
rect -155 2469 -36 2473
rect 76 2472 79 2476
rect 94 2472 114 2476
rect 246 2472 268 2476
rect 398 2472 422 2476
rect 550 2472 576 2476
rect 702 2472 730 2476
rect 854 2472 884 2476
rect 1006 2472 1038 2476
rect 1158 2472 1192 2476
rect 1310 2472 1346 2476
rect 1462 2472 1500 2476
rect 1614 2472 1654 2476
rect 1766 2472 1808 2476
rect 1918 2472 1962 2476
rect 2070 2472 2116 2476
rect 2222 2472 2270 2476
rect -155 2461 -36 2465
rect 76 2464 79 2468
rect 79 2457 83 2464
rect -155 2453 83 2457
rect 110 2427 114 2472
rect 264 2427 268 2472
rect 418 2427 422 2472
rect 572 2427 576 2472
rect 726 2427 730 2472
rect 880 2427 884 2472
rect 1034 2427 1038 2472
rect 1188 2427 1192 2472
rect 1342 2427 1346 2472
rect 1496 2427 1500 2472
rect 1650 2427 1654 2472
rect 1804 2427 1808 2472
rect 1958 2427 1962 2472
rect 2112 2427 2116 2472
rect 2266 2427 2270 2472
rect 2346 2455 2350 2480
rect 2354 2468 2358 2480
rect 2378 2481 2382 2488
rect 2406 2477 2427 2481
rect 2378 2476 2382 2477
rect 2366 2472 2382 2476
rect 2358 2464 2427 2468
rect 2346 2451 2427 2455
rect 2366 2438 2424 2442
rect 2420 2427 2424 2438
rect -148 2421 -125 2427
rect -155 2374 -36 2378
rect 2420 2374 2424 2378
rect -155 2359 -36 2363
rect -155 2351 -36 2355
rect 2434 2318 2437 2533
rect 2428 2315 2437 2318
rect 2440 2312 2443 2521
rect 2428 2309 2443 2312
rect 2446 2306 2449 2521
rect 2428 2303 2449 2306
rect 2452 2300 2455 2521
rect 2428 2297 2455 2300
rect 2458 2294 2461 2521
rect 2428 2291 2461 2294
rect 2464 2288 2467 2521
rect 2428 2285 2467 2288
rect 2470 2282 2473 2521
rect 2428 2279 2473 2282
rect 2476 2276 2479 2521
rect 2428 2273 2479 2276
rect 2482 2270 2485 2521
rect 2428 2267 2485 2270
rect 2488 2264 2491 2521
rect 2428 2261 2491 2264
rect 2494 2258 2497 2521
rect 2428 2255 2497 2258
rect 2500 2252 2503 2521
rect 2428 2249 2503 2252
rect 2506 2246 2509 2521
rect 2428 2243 2509 2246
rect 2512 2240 2515 2521
rect 2428 2237 2515 2240
rect 2518 2234 2521 2521
rect 2428 2231 2521 2234
rect 2524 2228 2527 2521
rect 2530 2481 2534 2521
rect 2534 2477 2568 2481
rect 2534 2464 2568 2468
rect 2541 2451 2568 2455
rect 2530 2355 2534 2451
rect 2541 2359 2568 2363
rect 2530 2351 2537 2355
rect 2541 2351 2568 2355
rect 2428 2225 2527 2228
use pin  pin_0
timestamp 1383821139
transform 1 0 413 0 1 2522
box -460 -103 2121 1847
use shift  shift_0
timestamp 1383822934
transform 1 0 154 0 1 2185
box -197 40 2282 342
<< labels >>
rlabel metal2 -155 2351 -147 2355 0 SCLKI
rlabel metal2 -155 2359 -147 2363 0 LDI
rlabel metal2 -155 2374 -147 2378 0 SI
rlabel metal2 -155 2469 -147 2473 0 PCLKI
rlabel metal2 -155 2461 -147 2465 0 PSI
rlabel metal2 2560 2351 2568 2355 0 SCLKO
rlabel metal2 2560 2359 2568 2363 0 LDO
rlabel metal2 2560 2581 2568 2585 0 PCLKO
rlabel metal2 2560 2477 2568 2481 0 PSO
rlabel metal2 2560 2464 2568 2468 0 TESTO
rlabel metal1 -139 2209 -131 2217 0 GND
rlabel metal1 -155 2193 -147 2201 0 VDD
rlabel metal2 2420 2374 2424 2378 0 SSO
rlabel metal2 -155 2453 -147 2457 0 TESTI
rlabel metal2 2560 2451 2568 2455 0 SO
<< end >>
