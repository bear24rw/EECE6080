magic
tech scmos
timestamp 1383903783
<< nwell >>
rect -12 4369 -11 4416
<< metal1 >>
rect -185 4481 2574 4491
rect -185 4367 -175 4481
rect -185 4361 -183 4367
rect -177 4361 -175 4367
rect -185 4251 -175 4361
rect -185 4245 -183 4251
rect -177 4245 -175 4251
rect -185 4135 -175 4245
rect -185 4129 -183 4135
rect -177 4129 -175 4135
rect -185 4019 -175 4129
rect -185 4013 -183 4019
rect -177 4013 -175 4019
rect -185 3903 -175 4013
rect -185 3897 -183 3903
rect -177 3897 -175 3903
rect -185 3787 -175 3897
rect -185 3781 -183 3787
rect -177 3781 -175 3787
rect -185 3671 -175 3781
rect -185 3665 -183 3671
rect -177 3665 -175 3671
rect -185 3555 -175 3665
rect -185 3549 -183 3555
rect -177 3549 -175 3555
rect -185 3439 -175 3549
rect -185 3433 -183 3439
rect -177 3433 -175 3439
rect -185 3323 -175 3433
rect -185 3317 -183 3323
rect -177 3317 -175 3323
rect -185 3207 -175 3317
rect -185 3201 -183 3207
rect -177 3201 -175 3207
rect -185 3091 -175 3201
rect -185 3085 -183 3091
rect -177 3085 -175 3091
rect -185 2975 -175 3085
rect -185 2969 -183 2975
rect -177 2969 -175 2975
rect -185 2859 -175 2969
rect -185 2853 -183 2859
rect -177 2853 -175 2859
rect -185 2743 -175 2853
rect -185 2737 -183 2743
rect -177 2737 -175 2743
rect -185 2627 -175 2737
rect -185 2621 -183 2627
rect -177 2621 -175 2627
rect -185 2427 -175 2621
rect -185 2421 -183 2427
rect -177 2421 -175 2427
rect -185 2194 -175 2421
rect -165 4461 2554 4471
rect -165 2214 -155 4461
rect -142 4361 -40 4367
rect 2544 4267 2554 4461
rect 2431 4261 2554 4267
rect -142 4245 -40 4251
rect 2544 4151 2554 4261
rect 2431 4145 2554 4151
rect -142 4129 -40 4135
rect 2544 4035 2554 4145
rect 2431 4029 2554 4035
rect -142 4013 -40 4019
rect 2544 3919 2554 4029
rect 2431 3913 2554 3919
rect -142 3897 -40 3903
rect 2544 3803 2554 3913
rect 2431 3797 2554 3803
rect -142 3781 -40 3787
rect 2544 3687 2554 3797
rect 2431 3681 2554 3687
rect -142 3665 -40 3671
rect 2544 3571 2554 3681
rect 2431 3565 2554 3571
rect -142 3549 -40 3555
rect 2544 3455 2554 3565
rect 2431 3449 2554 3455
rect -142 3433 -40 3439
rect 2544 3339 2554 3449
rect 2431 3333 2554 3339
rect -142 3317 -40 3323
rect 2544 3223 2554 3333
rect 2431 3217 2554 3223
rect -142 3201 -40 3207
rect 2544 3107 2554 3217
rect 2431 3101 2554 3107
rect -142 3085 -40 3091
rect 2544 2991 2554 3101
rect 2431 2985 2554 2991
rect -142 2969 -40 2975
rect 2544 2875 2554 2985
rect 2431 2869 2554 2875
rect -142 2853 -40 2859
rect 2544 2759 2554 2869
rect 2431 2753 2554 2759
rect -142 2737 -40 2743
rect 2544 2643 2554 2753
rect 2431 2637 2554 2643
rect -142 2621 -40 2627
rect 2432 2581 2537 2585
rect 2544 2527 2554 2637
rect 2431 2521 2554 2527
rect 2420 2487 2541 2491
rect 83 2480 2346 2484
rect 2358 2480 2374 2484
rect 2431 2477 2530 2481
rect 83 2472 2362 2476
rect 83 2464 2354 2468
rect 2362 2442 2366 2472
rect 2431 2464 2530 2468
rect 2537 2455 2541 2487
rect 2431 2451 2530 2455
rect -142 2421 -40 2427
rect 2431 2359 2537 2363
rect 2431 2351 2537 2355
rect 2544 2327 2554 2521
rect 2434 2321 2554 2327
rect -4 2221 0 2314
rect 150 2221 154 2314
rect 304 2221 308 2314
rect 458 2221 462 2314
rect 612 2221 616 2314
rect 1844 2221 1848 2314
rect 1998 2221 2002 2314
rect 2152 2221 2156 2314
rect 2306 2221 2310 2314
rect 2544 2214 2554 2321
rect -165 2204 2554 2214
rect 2564 2194 2574 4481
rect -185 2184 2574 2194
<< m2contact >>
rect -183 4361 -177 4367
rect -183 4245 -177 4251
rect -183 4129 -177 4135
rect -183 4013 -177 4019
rect -183 3897 -177 3903
rect -183 3781 -177 3787
rect -183 3665 -177 3671
rect -183 3549 -177 3555
rect -183 3433 -177 3439
rect -183 3317 -177 3323
rect -183 3201 -177 3207
rect -183 3085 -177 3091
rect -183 2969 -177 2975
rect -183 2853 -177 2859
rect -183 2737 -177 2743
rect -183 2621 -177 2627
rect -183 2421 -177 2427
rect -36 4437 -32 4441
rect -28 4427 -24 4431
rect 2415 4427 2419 4431
rect 2335 4417 2339 4421
rect 2391 4417 2395 4421
rect -148 4361 -142 4367
rect -148 4245 -142 4251
rect -148 4129 -142 4135
rect -148 4013 -142 4019
rect -148 3897 -142 3903
rect -148 3781 -142 3787
rect -148 3665 -142 3671
rect -148 3549 -142 3555
rect -148 3433 -142 3439
rect -148 3317 -142 3323
rect -148 3201 -142 3207
rect -148 3085 -142 3091
rect -148 2969 -142 2975
rect -148 2853 -142 2859
rect -148 2737 -142 2743
rect -148 2621 -142 2627
rect 2428 2581 2432 2585
rect 2537 2581 2541 2585
rect 79 2480 83 2484
rect 2346 2480 2350 2484
rect 2354 2480 2358 2484
rect 2378 2477 2382 2481
rect 2402 2477 2406 2481
rect 2427 2477 2431 2481
rect 2530 2477 2534 2481
rect 79 2472 83 2476
rect 2362 2472 2366 2476
rect 79 2464 83 2468
rect 2354 2464 2358 2468
rect 2427 2464 2431 2468
rect 2530 2464 2534 2468
rect 2427 2451 2431 2455
rect 2530 2451 2534 2455
rect 2537 2451 2541 2455
rect 2362 2438 2366 2442
rect -148 2421 -142 2427
rect 2427 2359 2431 2363
rect 2537 2359 2541 2363
rect 2427 2351 2431 2355
rect 2537 2351 2541 2355
rect -4 2217 0 2221
rect 150 2217 154 2221
rect 304 2217 308 2221
rect 458 2217 462 2221
rect 612 2217 616 2221
rect 1844 2217 1848 2221
rect 1998 2217 2002 2221
rect 2152 2217 2156 2221
rect 2306 2217 2310 2221
<< metal2 >>
rect -185 4437 -36 4441
rect -185 4427 -28 4431
rect -17 4387 -13 4491
rect -9 4407 -5 4491
rect -1 4451 3 4491
rect 94 4454 98 4491
rect 147 4455 151 4491
rect -9 4403 -1 4407
rect 155 4387 159 4491
rect 2149 4414 2153 4491
rect 2157 4429 2161 4491
rect 2165 4437 2169 4491
rect 2197 4467 2201 4491
rect 2157 4425 2165 4429
rect 2323 4414 2327 4491
rect 2335 4421 2339 4491
rect 2391 4421 2395 4491
rect 2415 4431 2419 4491
rect 2149 4410 2165 4414
rect 2319 4410 2327 4414
rect -17 4383 -1 4387
rect 151 4383 159 4387
rect -177 4361 -148 4367
rect -177 4245 -148 4251
rect -177 4129 -148 4135
rect -177 4013 -148 4019
rect -177 3897 -148 3903
rect -177 3781 -148 3787
rect -177 3665 -148 3671
rect -177 3549 -148 3555
rect -177 3433 -148 3439
rect -177 3317 -148 3323
rect -177 3201 -148 3207
rect -177 3085 -148 3091
rect -177 2969 -148 2975
rect -177 2853 -148 2859
rect -177 2737 -148 2743
rect -177 2621 -148 2627
rect 2541 2581 2574 2585
rect 2431 2533 2437 2537
rect 76 2480 79 2484
rect 94 2476 98 2530
rect 246 2476 250 2530
rect 398 2476 402 2530
rect 550 2476 554 2530
rect 702 2476 706 2530
rect 854 2476 858 2530
rect 1006 2476 1010 2530
rect 1158 2476 1162 2530
rect 1310 2476 1314 2530
rect 1462 2476 1466 2530
rect 1614 2476 1618 2530
rect 1766 2476 1770 2530
rect 1918 2476 1922 2530
rect 2070 2476 2074 2530
rect 2222 2476 2226 2530
rect 2374 2492 2378 2530
rect 2374 2488 2382 2492
rect -185 2469 -36 2473
rect 76 2472 79 2476
rect 94 2472 114 2476
rect 246 2472 268 2476
rect 398 2472 422 2476
rect 550 2472 576 2476
rect 702 2472 730 2476
rect 854 2472 884 2476
rect 1006 2472 1038 2476
rect 1158 2472 1192 2476
rect 1310 2472 1346 2476
rect 1462 2472 1500 2476
rect 1614 2472 1654 2476
rect 1766 2472 1808 2476
rect 1918 2472 1962 2476
rect 2070 2472 2116 2476
rect 2222 2472 2270 2476
rect -185 2461 -36 2465
rect 76 2464 79 2468
rect 79 2457 83 2464
rect -185 2453 83 2457
rect 110 2427 114 2472
rect 264 2427 268 2472
rect 418 2427 422 2472
rect 572 2427 576 2472
rect 726 2427 730 2472
rect 880 2427 884 2472
rect 1034 2427 1038 2472
rect 1188 2427 1192 2472
rect 1342 2427 1346 2472
rect 1496 2427 1500 2472
rect 1650 2427 1654 2472
rect 1804 2427 1808 2472
rect 1958 2427 1962 2472
rect 2112 2427 2116 2472
rect 2266 2427 2270 2472
rect 2346 2455 2350 2480
rect 2354 2468 2358 2480
rect 2378 2481 2382 2488
rect 2406 2477 2427 2481
rect 2378 2476 2382 2477
rect 2366 2472 2382 2476
rect 2358 2464 2427 2468
rect 2346 2451 2427 2455
rect 2366 2438 2424 2442
rect 2420 2427 2424 2438
rect -177 2421 -148 2427
rect -185 2374 -36 2378
rect 2420 2374 2424 2378
rect -185 2359 -36 2363
rect -185 2351 -36 2355
rect 2306 2318 2310 2319
rect 2434 2317 2437 2533
rect 2428 2314 2437 2317
rect 2440 2311 2443 2521
rect 2428 2308 2443 2311
rect 2446 2305 2449 2521
rect 2428 2302 2449 2305
rect 2452 2299 2455 2521
rect 2428 2296 2455 2299
rect 2458 2293 2461 2521
rect 2428 2290 2461 2293
rect 2464 2287 2467 2521
rect 2428 2284 2467 2287
rect 2470 2281 2473 2521
rect 2428 2278 2473 2281
rect 2476 2275 2479 2521
rect 2428 2272 2479 2275
rect 2482 2269 2485 2521
rect 2428 2266 2485 2269
rect 2488 2263 2491 2521
rect 2428 2260 2491 2263
rect 2494 2257 2497 2521
rect 2428 2254 2497 2257
rect 2500 2251 2503 2521
rect 2428 2248 2503 2251
rect 2506 2245 2509 2521
rect 2428 2242 2509 2245
rect 2512 2239 2515 2521
rect 2428 2236 2515 2239
rect 2518 2233 2521 2521
rect 2428 2230 2521 2233
rect 2524 2227 2527 2521
rect 2530 2481 2534 2521
rect 2534 2477 2574 2481
rect 2534 2464 2574 2468
rect 2541 2451 2574 2455
rect 2530 2355 2534 2451
rect 2541 2359 2574 2363
rect 2530 2351 2537 2355
rect 2541 2351 2574 2355
rect 2428 2224 2527 2227
rect -4 2184 0 2217
rect 150 2184 154 2217
rect 304 2184 308 2217
rect 458 2184 462 2217
rect 612 2184 616 2217
rect 1844 2184 1848 2217
rect 1998 2184 2002 2217
rect 2152 2184 2156 2217
rect 2306 2184 2310 2217
use INVX1_orig  INVX1_orig_0
timestamp 1053022145
transform 1 0 -38 0 -1 4464
box -9 -3 26 105
use pin_slice  pin_slice_0
timestamp 1383875311
transform 1 0 89 0 -1 4354
box -100 -113 68 -5
use shift_slice  shift_slice_0
timestamp 1383875311
transform 1 0 2174 0 -1 4467
box -16 0 151 108
use DFFPOSX1  DFFPOSX1_0
timestamp 1383875311
transform -1 0 2429 0 -1 4464
box -8 -3 104 105
use pin  pin_0
timestamp 1383882935
transform 1 0 413 0 1 2522
box -460 -103 2121 1847
use shift  shift_0
timestamp 1383882935
transform 1 0 154 0 1 2185
box -197 39 2282 342
<< labels >>
rlabel metal2 2420 2374 2424 2378 0 SSO
rlabel metal2 -185 2351 -175 2355 0 SCLKI
rlabel metal2 -185 2359 -175 2363 0 LDI
rlabel metal2 -185 2374 -175 2378 0 SI
rlabel metal2 -185 2453 -175 2457 0 TESTI
rlabel metal2 -185 2461 -175 2465 0 PSI
rlabel metal2 -185 2469 -175 2473 0 PCLKI
rlabel metal2 2564 2351 2574 2355 0 SCLKO
rlabel metal2 2564 2359 2574 2363 0 LDO
rlabel metal2 2564 2451 2574 2455 0 SO
rlabel metal2 2564 2464 2574 2468 0 TESTO
rlabel metal2 2564 2581 2574 2585 0 PCLKO
rlabel metal1 -165 2204 -155 2214 0 GND
rlabel metal1 -185 2184 -175 2194 0 VDD
rlabel metal2 -4 2184 0 2194 0 W0
rlabel metal2 150 2184 154 2194 0 W1
rlabel metal2 304 2184 308 2194 0 W2
rlabel metal2 458 2184 462 2194 0 W3
rlabel metal2 612 2184 616 2194 0 W4
rlabel metal2 1844 2184 1848 2194 0 W12
rlabel metal2 1998 2184 2002 2194 0 W13
rlabel metal2 2152 2184 2156 2194 0 W14
rlabel metal2 2306 2184 2310 2194 0 W15
rlabel metal2 -185 4437 -175 4441 0 TII
rlabel metal2 -185 4427 -175 4431 0 TIO
rlabel metal2 -17 4481 -13 4491 0 TPQI
rlabel metal2 -9 4481 -5 4491 0 TPCI
rlabel metal2 -1 4481 3 4491 0 TPZI
rlabel metal2 147 4481 151 4491 0 TPZO
rlabel metal2 155 4481 159 4491 0 TPQO
rlabel metal2 2149 4481 2153 4491 0 TSSI
rlabel metal2 2157 4481 2161 4491 0 TSLDI
rlabel metal2 2165 4481 2169 4491 0 TSCI
rlabel metal2 2197 4481 2201 4491 0 TSZ
rlabel metal2 2323 4481 2327 4491 0 TSSO
rlabel metal2 2335 4481 2339 4491 0 TFQ
rlabel metal2 2391 4481 2395 4491 0 TFD
rlabel metal2 2415 4481 2419 4491 0 TFC
rlabel metal2 94 4481 98 4491 0 TPWI
rlabel metal2 2564 2477 2574 2481 0 PSO
<< end >>
