magic
tech scmos
timestamp 1383634647
<< metal1 >>
rect -4 40 3 41
<< m2contact >>
rect -109 46 -105 50
rect -101 46 -97 50
rect -77 46 -73 50
rect -67 46 -63 50
rect -59 46 -55 50
rect -35 46 -31 50
rect -1 45 3 49
rect -77 36 -73 40
rect -35 36 -31 40
<< metal2 >>
rect -113 60 -55 64
rect -113 53 -97 57
rect -90 53 -63 57
rect -101 50 -97 53
rect -109 43 -105 46
rect -91 43 -87 53
rect -67 50 -63 53
rect -109 39 -87 43
rect -91 0 -87 39
rect -84 46 -77 50
rect -59 50 -55 60
rect -25 58 -21 1674
rect 2347 1670 2445 1674
rect 2347 1636 2438 1640
rect 2347 1520 2432 1524
rect 2347 1404 2426 1408
rect 2347 1288 2420 1292
rect 2347 1172 2414 1176
rect 2347 1056 2408 1060
rect 2347 940 2402 944
rect 2347 824 2396 828
rect 2347 708 2390 712
rect 2347 592 2384 596
rect 2347 476 2378 480
rect 2347 360 2372 364
rect 2347 244 2366 248
rect 2347 128 2360 132
rect -51 54 -21 58
rect -84 0 -80 46
rect -51 40 -47 54
rect -73 36 -47 40
rect -43 46 -35 50
rect -25 46 -21 54
rect -43 0 -39 46
rect -17 45 -1 49
rect -17 40 -13 45
rect -31 36 -13 40
rect 2347 37 2354 41
rect 2350 0 2354 37
rect 2357 0 2360 128
rect 2363 0 2366 244
rect 2369 0 2372 360
rect 2375 0 2378 476
rect 2381 0 2384 592
rect 2387 0 2390 708
rect 2393 0 2396 824
rect 2399 0 2402 940
rect 2405 0 2408 1056
rect 2411 0 2414 1172
rect 2417 0 2420 1288
rect 2423 0 2426 1404
rect 2429 0 2432 1520
rect 2435 0 2438 1636
rect 2441 0 2445 1670
use MUX2X1  MUX2X1_1
timestamp 1383629942
transform 1 0 -111 0 1 3
box -5 -3 53 105
use MUX2X1  MUX2X1_0
timestamp 1383629942
transform 1 0 -69 0 1 3
box -5 -3 53 105
use pin_buffer  pin_buffer_0
array 0 0 46 0 14 116
timestamp 1383629942
transform 1 0 -36 0 1 0
box 0 0 46 108
use pin_row_connect  pin_row_connect_0
array 0 0 98 0 13 116
timestamp 1383629942
transform 1 0 4 0 1 0
box -8 0 2347 165
use pin_slice  pin_slice_0
array 0 14 156 0 14 116
timestamp 1383629942
transform 1 0 100 0 1 113
box -100 -113 68 -5
<< labels >>
rlabel metal2 -113 60 -109 64 0 PSI
rlabel metal2 -113 53 -109 57 0 PCLKI
<< end >>
