magic
tech scmos
timestamp 1383810178
<< metal2 >>
rect -158 43 -154 136
rect -4 49 0 136
rect 150 55 154 136
rect 304 61 308 136
rect 458 67 462 136
rect 612 73 616 136
rect 766 79 770 136
rect 920 85 924 136
rect 1074 91 1078 136
rect 1228 97 1232 136
rect 1382 103 1386 136
rect 1536 109 1540 136
rect 1690 115 1694 136
rect 1844 121 1848 136
rect 1998 127 2002 136
rect 2152 133 2156 136
rect 2152 130 2274 133
rect 1998 124 2274 127
rect 1844 118 2274 121
rect 1690 112 2274 115
rect 1536 106 2274 109
rect 1382 100 2274 103
rect 1228 94 2274 97
rect 1074 88 2274 91
rect 920 82 2274 85
rect 766 76 2274 79
rect 612 70 2274 73
rect 458 64 2274 67
rect 304 58 2274 61
rect 150 52 2274 55
rect -4 46 2274 49
rect -158 40 2274 43
use mux  mux_0
timestamp 1383808422
transform 1 0 2209 0 -1 342
box 0 0 73 108
use shift_slice  shift_slice_0
array 0 15 154 0 0 108
timestamp 1383810178
transform 1 0 -181 0 1 136
box -16 0 151 108
<< end >>
