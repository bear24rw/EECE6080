magic
tech scmos
timestamp 1383808422
<< metal1 >>
rect 43 36 53 40
rect 49 30 53 36
use MUX2X1  MUX2X1_0
timestamp 1383808422
transform 1 0 5 0 1 3
box -5 -3 53 105
use INVX1  INVX1_0
timestamp 1383808422
transform 1 0 47 0 1 3
box -9 -3 26 105
<< end >>
