magic
tech scmos
timestamp 1383634647
<< nwell >>
rect -60 1839 -53 1845
rect -60 1723 -53 1729
rect -60 1607 -53 1613
rect -60 1491 -53 1497
rect -60 1375 -53 1381
rect -60 1259 -53 1265
rect -60 1143 -53 1149
rect -60 1027 -53 1033
rect -60 911 -53 917
rect -60 795 -53 801
rect -60 679 -53 685
rect -60 563 -53 569
rect -60 447 -53 453
<< metal1 >>
rect -171 1861 2445 1869
rect -171 1845 -163 1861
rect -171 1839 -170 1845
rect -164 1839 -163 1845
rect -171 1729 -163 1839
rect -171 1723 -170 1729
rect -164 1723 -163 1729
rect -171 1613 -163 1723
rect -171 1607 -170 1613
rect -164 1607 -163 1613
rect -171 1497 -163 1607
rect -171 1491 -170 1497
rect -164 1491 -163 1497
rect -171 1381 -163 1491
rect -171 1375 -170 1381
rect -164 1375 -163 1381
rect -171 1265 -163 1375
rect -171 1259 -170 1265
rect -164 1259 -163 1265
rect -171 1149 -163 1259
rect -171 1143 -170 1149
rect -164 1143 -163 1149
rect -171 1033 -163 1143
rect -171 1027 -170 1033
rect -164 1027 -163 1033
rect -171 917 -163 1027
rect -171 911 -170 917
rect -164 911 -163 917
rect -171 801 -163 911
rect -171 795 -170 801
rect -164 795 -163 801
rect -171 685 -163 795
rect -171 679 -170 685
rect -164 679 -163 685
rect -171 569 -163 679
rect -171 563 -170 569
rect -164 563 -163 569
rect -171 453 -163 563
rect -171 447 -170 453
rect -164 447 -163 453
rect -171 337 -163 447
rect -171 331 -170 337
rect -164 331 -163 337
rect -171 221 -163 331
rect -171 215 -170 221
rect -164 215 -163 221
rect -171 91 -163 215
rect -171 85 -170 91
rect -164 85 -163 91
rect -171 -121 -163 85
rect -159 1849 2433 1857
rect -159 -109 -151 1849
rect -142 1839 -53 1845
rect 2425 1745 2433 1849
rect 2322 1739 2433 1745
rect -142 1723 -53 1729
rect 2425 1629 2433 1739
rect 2322 1623 2433 1629
rect -142 1607 -53 1613
rect 2425 1513 2433 1623
rect 2322 1507 2433 1513
rect -142 1491 -53 1497
rect 2425 1397 2433 1507
rect 2322 1391 2433 1397
rect -142 1375 -53 1381
rect 2425 1281 2433 1391
rect 2322 1275 2433 1281
rect -142 1259 -53 1265
rect 2425 1165 2433 1275
rect 2322 1159 2433 1165
rect -142 1143 -53 1149
rect 2425 1049 2433 1159
rect 2322 1043 2433 1049
rect -142 1027 -53 1033
rect 2425 933 2433 1043
rect 2322 927 2433 933
rect -142 911 -53 917
rect 2425 817 2433 927
rect 2322 811 2433 817
rect -142 795 -53 801
rect 2425 701 2433 811
rect 2322 695 2433 701
rect -142 679 -53 685
rect 2425 585 2433 695
rect 2322 579 2433 585
rect -142 563 -53 569
rect 2425 469 2433 579
rect 2322 463 2433 469
rect -142 447 -53 453
rect 2425 353 2433 463
rect 2322 347 2433 353
rect -142 331 -53 337
rect 2425 237 2433 347
rect 2322 231 2433 237
rect -142 215 -137 221
rect 2425 121 2433 231
rect 2320 115 2433 121
rect -63 108 2288 112
rect 2310 108 2417 112
rect -104 101 2281 105
rect 2285 101 2417 105
rect -111 94 2295 98
rect 2299 94 2417 98
rect 2330 87 2417 91
rect 2317 28 2417 32
rect 2310 21 2417 25
rect 2425 -9 2433 115
rect 2320 -15 2433 -9
rect 2425 -109 2433 -15
rect -159 -117 2433 -109
rect 2437 -121 2445 1861
rect -171 -129 2445 -121
<< m2contact >>
rect -170 1839 -164 1845
rect -170 1723 -164 1729
rect -170 1607 -164 1613
rect -170 1491 -164 1497
rect -170 1375 -164 1381
rect -170 1259 -164 1265
rect -170 1143 -164 1149
rect -170 1027 -164 1033
rect -170 911 -164 917
rect -170 795 -164 801
rect -170 679 -164 685
rect -170 563 -164 569
rect -170 447 -164 453
rect -170 331 -164 337
rect -170 215 -164 221
rect -170 85 -164 91
rect -148 1839 -142 1845
rect -148 1723 -142 1729
rect -148 1607 -142 1613
rect -148 1491 -142 1497
rect -148 1375 -142 1381
rect -148 1259 -142 1265
rect -148 1143 -142 1149
rect -148 1027 -142 1033
rect -148 911 -142 917
rect -148 795 -142 801
rect -148 679 -142 685
rect -148 563 -142 569
rect -148 447 -142 453
rect -148 331 -142 337
rect -148 215 -142 221
rect -67 108 -63 112
rect 2288 108 2292 112
rect 2306 108 2310 112
rect 2417 108 2421 112
rect -108 101 -104 105
rect 2281 101 2285 105
rect 2417 101 2421 105
rect -115 94 -111 98
rect 2295 94 2299 98
rect 2417 94 2421 98
rect -148 85 -142 91
rect 2326 87 2330 91
rect 2417 87 2421 91
rect 2306 31 2310 35
rect 2313 28 2317 32
rect 2417 28 2421 32
rect 2417 21 2421 25
<< metal2 >>
rect -164 1839 -148 1845
rect -164 1723 -148 1729
rect -164 1607 -148 1613
rect -164 1491 -148 1497
rect -164 1375 -148 1381
rect -164 1259 -148 1265
rect -164 1143 -148 1149
rect -164 1027 -148 1033
rect -164 911 -148 917
rect -164 795 -148 801
rect -164 679 -148 685
rect -164 563 -148 569
rect -164 447 -148 453
rect -164 331 -148 337
rect -164 215 -148 221
rect -171 175 -137 179
rect -171 168 -137 172
rect -115 98 -111 115
rect -108 105 -104 115
rect -67 112 -63 115
rect 81 105 85 124
rect 237 105 241 124
rect 393 105 397 124
rect 549 105 553 124
rect 705 105 709 124
rect 861 105 865 124
rect 1017 105 1021 124
rect 1173 105 1177 124
rect 1329 105 1333 124
rect 1485 105 1489 124
rect 1641 105 1645 124
rect 1797 105 1801 124
rect 1953 105 1957 124
rect 2109 105 2113 124
rect 13 101 85 105
rect 174 101 241 105
rect 335 101 397 105
rect 496 101 553 105
rect 657 101 709 105
rect 818 101 865 105
rect 979 101 1021 105
rect 1140 101 1177 105
rect 1301 101 1333 105
rect 1462 101 1489 105
rect 1623 101 1645 105
rect 1784 101 1801 105
rect 1945 101 1957 105
rect 2106 101 2113 105
rect 2265 105 2269 128
rect 2274 115 2317 119
rect 2265 101 2271 105
rect -171 94 -115 98
rect 13 91 17 101
rect 174 91 178 101
rect 335 91 339 101
rect 496 91 500 101
rect 657 91 661 101
rect 818 91 822 101
rect 979 91 983 101
rect 1140 91 1144 101
rect 1301 91 1305 101
rect 1462 91 1466 101
rect 1623 91 1627 101
rect 1784 91 1788 101
rect 1945 91 1949 101
rect 2106 91 2110 101
rect 2267 91 2271 101
rect 2274 91 2278 115
rect 2281 91 2285 101
rect 2288 91 2292 108
rect 2295 91 2299 94
rect -164 85 -148 91
rect -171 71 -145 75
rect -171 64 -145 68
rect -171 38 -145 42
rect 2306 35 2310 108
rect 2313 32 2317 115
rect 2320 -18 2323 127
rect 2326 91 2330 115
rect 2312 -21 2323 -18
rect 2333 -24 2336 115
rect 2312 -27 2336 -24
rect 2339 -30 2342 115
rect 2312 -33 2342 -30
rect 2345 -36 2348 115
rect 2312 -39 2348 -36
rect 2351 -42 2354 115
rect 2312 -45 2354 -42
rect 2357 -48 2360 115
rect 2312 -51 2360 -48
rect 2363 -54 2366 115
rect 2312 -57 2366 -54
rect 2369 -60 2372 115
rect 2312 -63 2372 -60
rect 2375 -66 2378 115
rect 2312 -69 2378 -66
rect 2381 -72 2384 115
rect 2312 -75 2384 -72
rect 2387 -78 2390 115
rect 2312 -81 2390 -78
rect 2393 -84 2396 115
rect 2312 -87 2396 -84
rect 2399 -90 2402 115
rect 2312 -93 2402 -90
rect 2405 -96 2408 115
rect 2312 -99 2408 -96
rect 2411 -102 2414 115
rect 2417 112 2421 115
rect 2421 108 2445 112
rect 2421 101 2445 105
rect 2421 94 2445 98
rect 2421 87 2445 91
rect 2421 28 2445 32
rect 2421 21 2445 25
rect 2312 -105 2414 -102
use pin  pin_0
timestamp 1383634647
transform 1 0 -24 0 1 115
box -116 0 2445 1732
use shift  shift_0
timestamp 1383634647
transform 1 0 -128 0 1 -19
box -17 -86 2453 112
<< labels >>
rlabel metal2 -171 168 -163 172 0 PCLKI
rlabel metal2 -171 175 -163 179 0 PSI
rlabel metal2 -171 71 -163 75 0 LDI
rlabel metal2 -171 64 -163 68 0 SCLKI
rlabel metal2 -171 38 -163 42 0 SI
rlabel metal2 -171 94 -163 98 0 TESTI
rlabel metal2 2437 108 2445 112 0 PSO
rlabel metal2 2437 21 2445 25 0 SO
rlabel metal2 2437 94 2445 98 0 TESTO
rlabel metal2 2437 101 2445 105 0 SCLKO
rlabel metal2 2437 28 2445 32 0 LDO
rlabel metal2 2437 87 2445 91 0 PCLKO
<< end >>
