magic
tech scmos
timestamp 1383634647
use top  top_0
timestamp 1383634647
transform 1 0 1364 0 1 1679
box -171 -129 2445 1869
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1072203966
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< end >>
