magic
tech scmos
timestamp 1383792416
<< nwell >>
rect -60 1839 -53 1845
rect -60 1723 -53 1729
rect -60 1607 -53 1613
rect -60 1491 -53 1497
rect -60 1375 -53 1381
rect -60 1259 -53 1265
rect -60 1143 -53 1149
rect -60 1027 -53 1033
rect -60 911 -53 917
rect -60 795 -53 801
rect -60 679 -53 685
rect -60 563 -53 569
rect -60 447 -53 453
<< metal1 >>
rect -198 1861 2445 1869
rect -198 1845 -190 1861
rect -198 1839 -197 1845
rect -191 1839 -190 1845
rect -198 1729 -190 1839
rect -198 1723 -197 1729
rect -191 1723 -190 1729
rect -198 1613 -190 1723
rect -198 1607 -197 1613
rect -191 1607 -190 1613
rect -198 1497 -190 1607
rect -198 1491 -197 1497
rect -191 1491 -190 1497
rect -198 1381 -190 1491
rect -198 1375 -197 1381
rect -191 1375 -190 1381
rect -198 1265 -190 1375
rect -198 1259 -197 1265
rect -191 1259 -190 1265
rect -198 1149 -190 1259
rect -198 1143 -197 1149
rect -191 1143 -190 1149
rect -198 1033 -190 1143
rect -198 1027 -197 1033
rect -191 1027 -190 1033
rect -198 917 -190 1027
rect -198 911 -197 917
rect -191 911 -190 917
rect -198 801 -190 911
rect -198 795 -197 801
rect -191 795 -190 801
rect -198 685 -190 795
rect -198 679 -197 685
rect -191 679 -190 685
rect -198 569 -190 679
rect -198 563 -197 569
rect -191 563 -190 569
rect -198 453 -190 563
rect -198 447 -197 453
rect -191 447 -190 453
rect -198 337 -190 447
rect -198 331 -197 337
rect -191 331 -190 337
rect -198 221 -190 331
rect -198 215 -197 221
rect -191 215 -190 221
rect -198 91 -190 215
rect -198 85 -197 91
rect -191 85 -190 91
rect -198 -121 -190 85
rect -186 1849 2433 1857
rect -186 -109 -178 1849
rect -169 1839 -53 1845
rect 2425 1745 2433 1849
rect 2322 1739 2433 1745
rect -169 1723 -53 1729
rect 2425 1629 2433 1739
rect 2322 1623 2433 1629
rect -169 1607 -53 1613
rect 2425 1513 2433 1623
rect 2322 1507 2433 1513
rect -169 1491 -53 1497
rect 2425 1397 2433 1507
rect 2322 1391 2433 1397
rect -169 1375 -53 1381
rect 2425 1281 2433 1391
rect 2322 1275 2433 1281
rect -169 1259 -53 1265
rect 2425 1165 2433 1275
rect 2322 1159 2433 1165
rect -169 1143 -53 1149
rect 2425 1049 2433 1159
rect 2322 1043 2433 1049
rect -169 1027 -53 1033
rect 2425 933 2433 1043
rect 2322 927 2433 933
rect -169 911 -53 917
rect 2425 817 2433 927
rect 2322 811 2433 817
rect -169 795 -53 801
rect 2425 701 2433 811
rect 2322 695 2433 701
rect -169 679 -53 685
rect 2425 585 2433 695
rect 2322 579 2433 585
rect -169 563 -53 569
rect 2425 469 2433 579
rect 2322 463 2433 469
rect -169 447 -53 453
rect 2425 353 2433 463
rect 2322 347 2433 353
rect -169 331 -53 337
rect 2425 237 2433 347
rect 2322 231 2433 237
rect 2425 121 2433 231
rect 2320 115 2433 121
rect -71 108 2292 112
rect 2310 108 2417 112
rect -129 101 2285 105
rect 2289 101 2417 105
rect -145 94 2299 98
rect 2303 94 2417 98
rect 2330 87 2417 91
rect 2317 80 2417 84
rect 2313 73 2417 77
rect 2313 25 2317 73
rect 2304 21 2317 25
rect 2425 -9 2433 115
rect 2308 -15 2433 -9
rect 2425 -109 2433 -15
rect -186 -117 2433 -109
rect 2437 -121 2445 1861
rect -198 -129 2445 -121
<< m2contact >>
rect -197 1839 -191 1845
rect -197 1723 -191 1729
rect -197 1607 -191 1613
rect -197 1491 -191 1497
rect -197 1375 -191 1381
rect -197 1259 -191 1265
rect -197 1143 -191 1149
rect -197 1027 -191 1033
rect -197 911 -191 917
rect -197 795 -191 801
rect -197 679 -191 685
rect -197 563 -191 569
rect -197 447 -191 453
rect -197 331 -191 337
rect -197 215 -191 221
rect -197 85 -191 91
rect -175 1839 -169 1845
rect -175 1723 -169 1729
rect -175 1607 -169 1613
rect -175 1491 -169 1497
rect -175 1375 -169 1381
rect -175 1259 -169 1265
rect -175 1143 -169 1149
rect -175 1027 -169 1033
rect -175 911 -169 917
rect -175 795 -169 801
rect -175 679 -169 685
rect -175 563 -169 569
rect -175 447 -169 453
rect -175 331 -169 337
rect -175 215 -169 221
rect -75 108 -71 112
rect 2292 108 2296 112
rect 2306 108 2310 112
rect 2417 108 2421 112
rect -133 101 -129 105
rect 2285 101 2289 105
rect 2417 101 2421 105
rect -149 94 -145 98
rect 2299 94 2303 98
rect 2417 94 2421 98
rect -175 85 -169 91
rect 2326 87 2330 91
rect 2417 87 2421 91
rect 2313 80 2317 84
rect 2417 80 2421 84
rect 2417 73 2421 77
rect 2282 31 2286 35
<< metal2 >>
rect -191 1839 -175 1845
rect -191 1723 -175 1729
rect -191 1607 -175 1613
rect -191 1491 -175 1497
rect -191 1375 -175 1381
rect -191 1259 -175 1265
rect -191 1143 -175 1149
rect -191 1027 -175 1033
rect -191 911 -175 917
rect -191 795 -175 801
rect -191 679 -175 685
rect -191 563 -175 569
rect -191 447 -175 453
rect -191 331 -175 337
rect -191 215 -175 221
rect -198 175 -169 179
rect -198 168 -169 172
rect -149 98 -145 115
rect -133 105 -129 115
rect -75 112 -71 115
rect 81 105 85 124
rect 237 105 241 124
rect 393 105 397 124
rect 549 105 553 124
rect 705 105 709 124
rect 861 105 865 124
rect 1017 105 1021 124
rect 1173 105 1177 124
rect 1329 105 1333 124
rect 1485 105 1489 124
rect 1641 105 1645 124
rect 1797 105 1801 124
rect 1953 105 1957 124
rect 2109 105 2113 124
rect 2265 105 2269 128
rect -11 101 85 105
rect 150 101 241 105
rect 311 101 397 105
rect 472 101 553 105
rect 633 101 709 105
rect 794 101 865 105
rect 955 101 1021 105
rect 1116 101 1177 105
rect 1277 101 1333 105
rect 1438 101 1489 105
rect 1599 101 1645 105
rect 1760 101 1801 105
rect 1921 101 1957 105
rect 2082 101 2113 105
rect 2243 101 2269 105
rect 2278 115 2317 119
rect -198 94 -149 98
rect -11 91 -7 101
rect 150 91 154 101
rect 311 91 315 101
rect 472 91 476 101
rect 633 91 637 101
rect 794 91 798 101
rect 955 91 959 101
rect 1116 91 1120 101
rect 1277 91 1281 101
rect 1438 91 1442 101
rect 1599 91 1603 101
rect 1760 91 1764 101
rect 1921 91 1925 101
rect 2082 91 2086 101
rect 2243 91 2247 101
rect 2278 91 2282 115
rect 2285 91 2289 101
rect 2292 91 2296 108
rect 2299 91 2303 94
rect -191 85 -175 91
rect -198 71 -169 75
rect -198 64 -169 68
rect -198 38 -169 42
rect 2243 38 2253 42
rect 2306 35 2310 108
rect 2313 84 2317 115
rect 2286 31 2310 35
rect 2320 -18 2323 127
rect 2326 91 2330 115
rect 2316 -21 2323 -18
rect 2333 -24 2336 115
rect 2316 -27 2336 -24
rect 2339 -30 2342 115
rect 2316 -33 2342 -30
rect 2345 -36 2348 115
rect 2316 -39 2348 -36
rect 2351 -42 2354 115
rect 2316 -45 2354 -42
rect 2357 -48 2360 115
rect 2316 -51 2360 -48
rect 2363 -54 2366 115
rect 2316 -57 2366 -54
rect 2369 -60 2372 115
rect 2316 -63 2372 -60
rect 2375 -66 2378 115
rect 2316 -69 2378 -66
rect 2381 -72 2384 115
rect 2316 -75 2384 -72
rect 2387 -78 2390 115
rect 2316 -81 2390 -78
rect 2393 -84 2396 115
rect 2316 -87 2396 -84
rect 2399 -90 2402 115
rect 2316 -93 2402 -90
rect 2405 -96 2408 115
rect 2316 -99 2408 -96
rect 2411 -102 2414 115
rect 2417 112 2421 115
rect 2421 108 2445 112
rect 2421 101 2445 105
rect 2421 94 2445 98
rect 2421 87 2445 91
rect 2421 80 2445 84
rect 2421 73 2445 77
rect 2316 -105 2414 -102
use pin  pin_0
timestamp 1383792416
transform 1 0 -24 0 1 115
box -148 0 2445 1732
use shift  shift_0
timestamp 1383647326
transform 1 0 -152 0 1 -19
box -17 -86 2468 112
<< labels >>
rlabel metal2 2437 108 2445 112 0 PSO
rlabel metal2 2437 94 2445 98 0 TESTO
rlabel metal2 2437 101 2445 105 0 SCLKO
rlabel metal2 2437 87 2445 91 0 PCLKO
rlabel metal2 2437 80 2445 84 0 LDO
rlabel metal2 2437 73 2445 77 0 SO
rlabel metal1 -186 -117 -178 -109 0 GND
rlabel metal1 -198 -129 -190 -121 0 VDD
rlabel metal2 -198 94 -190 98 0 TESTI
rlabel metal2 -198 38 -190 42 0 SI
rlabel metal2 -198 64 -190 68 0 SCLKI
rlabel metal2 -198 71 -190 75 0 LDI
rlabel metal2 -198 175 -190 179 0 PSI
rlabel metal2 -198 168 -190 172 0 PCLKI
rlabel metal2 2243 38 2253 42 0 SSO
<< end >>
