magic
tech scmos
timestamp 1383829970
<< metal1 >>
rect 15 147 435 189
rect 15 78 36 147
rect 57 146 77 147
rect 57 145 76 146
rect 57 144 75 145
rect 57 143 74 144
rect 57 142 73 143
rect 57 141 72 142
rect 57 140 71 141
rect 57 139 70 140
rect 57 138 69 139
rect 57 137 68 138
rect 57 136 67 137
rect 57 135 66 136
rect 57 78 63 135
rect 108 129 114 147
rect 159 129 165 147
rect 199 146 231 147
rect 200 145 231 146
rect 201 144 231 145
rect 264 144 279 147
rect 202 143 228 144
rect 203 142 228 143
rect 204 141 228 142
rect 264 141 276 144
rect 205 140 225 141
rect 206 139 225 140
rect 207 138 225 139
rect 208 137 225 138
rect 209 136 225 137
rect 210 135 225 136
rect 264 138 273 141
rect 264 135 270 138
rect 211 134 222 135
rect 212 133 222 134
rect 213 132 222 133
rect 264 132 267 135
rect 84 78 90 129
rect 108 117 126 129
rect 111 78 126 117
rect 15 69 126 78
rect 147 78 165 129
rect 186 117 192 129
rect 213 126 219 132
rect 213 123 216 126
rect 240 123 243 129
rect 210 111 216 123
rect 237 120 243 123
rect 198 108 216 111
rect 204 105 216 108
rect 186 99 189 105
rect 207 102 216 105
rect 186 78 192 99
rect 147 69 192 78
rect 210 78 216 102
rect 237 78 243 108
rect 261 78 267 132
rect 288 78 294 129
rect 312 78 318 147
rect 363 129 369 147
rect 336 117 369 129
rect 390 120 396 147
rect 417 120 435 147
rect 414 117 435 120
rect 348 108 369 117
rect 411 114 435 117
rect 405 111 435 114
rect 405 108 408 111
rect 348 105 381 108
rect 336 102 378 105
rect 336 99 375 102
rect 336 96 372 99
rect 336 93 369 96
rect 363 78 369 93
rect 390 78 396 99
rect 417 78 435 111
rect 210 69 435 78
rect 15 18 435 69
<< metal2 >>
rect 0 189 450 204
rect 0 183 18 189
rect 51 186 60 189
rect 93 186 102 189
rect 48 183 63 186
rect 90 183 105 186
rect 135 183 147 189
rect 177 183 189 189
rect 219 183 231 189
rect 261 183 273 189
rect 303 183 315 189
rect 348 186 357 189
rect 390 186 399 189
rect 345 183 360 186
rect 387 183 402 186
rect 432 183 450 189
rect 0 180 21 183
rect 45 180 54 183
rect 57 180 66 183
rect 87 180 96 183
rect 99 180 108 183
rect 132 180 150 183
rect 174 180 192 183
rect 216 180 234 183
rect 258 180 276 183
rect 300 180 318 183
rect 342 180 363 183
rect 384 180 405 183
rect 429 180 450 183
rect 0 153 15 180
rect 18 177 24 180
rect 42 177 51 180
rect 60 177 69 180
rect 84 177 93 180
rect 102 177 111 180
rect 129 177 135 180
rect 144 177 153 180
rect 171 177 177 180
rect 186 177 195 180
rect 213 177 222 180
rect 228 177 237 180
rect 255 177 264 180
rect 273 177 279 180
rect 297 177 306 180
rect 315 177 321 180
rect 339 177 348 180
rect 357 177 366 180
rect 381 177 390 180
rect 399 177 408 180
rect 426 177 432 180
rect 21 174 27 177
rect 39 174 48 177
rect 63 174 72 177
rect 81 174 90 177
rect 105 174 114 177
rect 126 174 132 177
rect 147 174 156 177
rect 168 174 174 177
rect 189 174 198 177
rect 210 174 219 177
rect 231 174 240 177
rect 252 174 261 177
rect 276 174 282 177
rect 294 174 303 177
rect 318 174 324 177
rect 336 174 345 177
rect 360 174 369 177
rect 378 174 387 177
rect 402 174 411 177
rect 423 174 429 177
rect 24 171 30 174
rect 36 171 45 174
rect 66 171 75 174
rect 78 171 87 174
rect 108 171 117 174
rect 123 171 129 174
rect 150 171 159 174
rect 165 171 171 174
rect 192 171 201 174
rect 207 171 216 174
rect 234 171 243 174
rect 249 171 258 174
rect 279 171 285 174
rect 291 171 300 174
rect 321 171 327 174
rect 333 171 342 174
rect 363 171 372 174
rect 375 171 384 174
rect 405 171 414 174
rect 420 171 426 174
rect 27 168 42 171
rect 69 168 84 171
rect 111 168 126 171
rect 153 168 168 171
rect 195 168 213 171
rect 237 168 255 171
rect 282 168 297 171
rect 324 168 339 171
rect 366 168 381 171
rect 408 168 423 171
rect 30 165 39 168
rect 72 165 81 168
rect 114 165 123 168
rect 27 162 39 165
rect 69 162 84 165
rect 114 162 126 165
rect 156 162 168 168
rect 198 162 210 168
rect 240 162 252 168
rect 282 162 294 168
rect 327 165 336 168
rect 369 165 378 168
rect 411 165 420 168
rect 324 162 336 165
rect 366 162 381 165
rect 411 162 423 165
rect 24 159 42 162
rect 66 159 87 162
rect 111 159 129 162
rect 153 159 171 162
rect 195 159 213 162
rect 237 159 255 162
rect 279 159 297 162
rect 321 159 339 162
rect 363 159 384 162
rect 408 159 426 162
rect 21 156 30 159
rect 39 156 45 159
rect 63 156 72 159
rect 81 156 90 159
rect 108 156 114 159
rect 123 156 132 159
rect 150 156 156 159
rect 165 156 174 159
rect 192 156 201 159
rect 207 156 216 159
rect 234 156 243 159
rect 249 156 258 159
rect 276 156 285 159
rect 294 156 300 159
rect 318 156 327 159
rect 336 156 342 159
rect 360 156 369 159
rect 378 156 387 159
rect 405 156 411 159
rect 420 156 429 159
rect 18 153 27 156
rect 42 153 48 156
rect 60 153 69 156
rect 84 153 93 156
rect 105 153 111 156
rect 126 153 135 156
rect 147 153 153 156
rect 168 153 177 156
rect 189 153 198 156
rect 210 153 219 156
rect 231 153 240 156
rect 252 153 261 156
rect 273 153 282 156
rect 297 153 303 156
rect 315 153 324 156
rect 339 153 345 156
rect 357 153 366 156
rect 381 153 390 156
rect 402 153 408 156
rect 423 153 432 156
rect 435 153 450 180
rect 0 150 24 153
rect 45 150 51 153
rect 57 150 66 153
rect 87 150 96 153
rect 102 150 108 153
rect 129 150 138 153
rect 144 150 150 153
rect 171 150 180 153
rect 186 150 195 153
rect 213 150 222 153
rect 228 150 237 153
rect 255 150 264 153
rect 270 150 279 153
rect 300 150 306 153
rect 312 150 321 153
rect 342 150 348 153
rect 354 150 363 153
rect 384 150 393 153
rect 399 150 405 153
rect 426 150 450 153
rect 0 147 21 150
rect 33 147 63 150
rect 74 149 202 150
rect 73 148 203 149
rect 72 147 204 148
rect 216 147 420 150
rect 429 147 450 150
rect 0 141 18 147
rect 0 138 21 141
rect 0 111 15 138
rect 18 135 24 138
rect 21 132 27 135
rect 30 132 36 147
rect 24 129 36 132
rect 27 126 36 129
rect 30 123 36 126
rect 27 120 36 123
rect 24 117 36 120
rect 21 114 36 117
rect 18 111 27 114
rect 0 108 24 111
rect 0 105 21 108
rect 0 99 18 105
rect 0 96 21 99
rect 0 93 24 96
rect 0 66 15 93
rect 18 90 27 93
rect 30 90 36 114
rect 21 87 36 90
rect 24 84 36 87
rect 27 81 36 84
rect 30 78 36 81
rect 57 141 60 147
rect 71 146 77 147
rect 70 145 76 146
rect 69 144 75 145
rect 68 143 74 144
rect 67 142 73 143
rect 66 141 72 142
rect 57 140 71 141
rect 57 139 70 140
rect 57 138 69 139
rect 57 137 68 138
rect 57 136 67 137
rect 57 135 66 136
rect 57 78 63 135
rect 108 129 114 147
rect 159 129 165 147
rect 199 146 205 147
rect 200 145 206 146
rect 201 144 207 145
rect 219 144 231 147
rect 264 144 279 147
rect 202 143 208 144
rect 203 142 209 143
rect 204 141 210 142
rect 219 141 228 144
rect 264 141 276 144
rect 205 140 211 141
rect 206 139 212 140
rect 207 138 213 139
rect 216 138 225 141
rect 208 137 225 138
rect 209 136 225 137
rect 210 135 225 136
rect 264 138 273 141
rect 264 135 270 138
rect 211 134 222 135
rect 212 133 222 134
rect 213 132 222 133
rect 264 132 267 135
rect 84 78 90 129
rect 108 117 126 129
rect 111 87 114 117
rect 120 87 126 117
rect 111 78 126 87
rect 27 75 126 78
rect 24 72 117 75
rect 21 69 27 72
rect 30 69 114 72
rect 120 69 126 75
rect 147 114 165 129
rect 186 117 192 129
rect 213 126 219 132
rect 213 123 216 126
rect 240 123 243 129
rect 147 111 156 114
rect 147 108 153 111
rect 147 96 150 108
rect 147 93 153 96
rect 147 90 156 93
rect 159 90 165 114
rect 210 111 216 123
rect 237 120 243 123
rect 198 108 216 111
rect 204 105 216 108
rect 147 87 165 90
rect 147 75 150 87
rect 153 84 165 87
rect 156 78 165 84
rect 186 99 189 105
rect 207 102 216 105
rect 186 78 192 99
rect 153 75 192 78
rect 147 72 192 75
rect 147 69 156 72
rect 159 69 192 72
rect 210 78 216 102
rect 237 78 243 105
rect 261 78 267 132
rect 288 78 294 129
rect 312 78 318 147
rect 363 129 369 147
rect 336 117 369 129
rect 390 120 396 147
rect 417 132 420 147
rect 432 141 450 147
rect 429 138 450 141
rect 426 135 432 138
rect 423 132 429 135
rect 417 129 426 132
rect 417 120 423 129
rect 414 117 426 120
rect 348 108 351 117
rect 363 114 369 117
rect 411 114 429 117
rect 360 111 369 114
rect 357 108 369 111
rect 405 111 420 114
rect 423 111 432 114
rect 435 111 450 138
rect 405 108 408 111
rect 348 105 360 108
rect 363 105 369 108
rect 336 99 357 105
rect 363 102 378 105
rect 363 99 375 102
rect 336 96 360 99
rect 363 96 372 99
rect 336 93 369 96
rect 363 78 369 93
rect 390 78 396 99
rect 417 90 420 111
rect 426 108 450 111
rect 429 105 450 108
rect 432 99 450 105
rect 429 96 450 99
rect 426 93 450 96
rect 423 90 432 93
rect 417 87 429 90
rect 417 84 426 87
rect 417 78 423 84
rect 210 75 423 78
rect 210 72 426 75
rect 210 69 420 72
rect 423 69 429 72
rect 18 66 24 69
rect 30 66 111 69
rect 120 66 153 69
rect 159 66 417 69
rect 426 66 432 69
rect 435 66 450 93
rect 0 63 21 66
rect 45 63 63 66
rect 90 63 108 66
rect 0 57 18 63
rect 48 60 60 63
rect 51 57 60 60
rect 93 60 105 63
rect 120 60 150 66
rect 174 63 234 66
rect 258 63 276 66
rect 300 63 318 66
rect 342 63 360 66
rect 387 63 405 66
rect 429 63 450 66
rect 177 60 216 63
rect 93 57 102 60
rect 120 57 147 60
rect 177 57 213 60
rect 219 57 231 63
rect 261 57 273 63
rect 303 57 315 63
rect 345 60 357 63
rect 348 57 357 60
rect 390 60 402 63
rect 390 57 399 60
rect 432 57 450 63
rect 0 54 21 57
rect 48 54 63 57
rect 90 54 105 57
rect 132 54 147 57
rect 174 54 192 57
rect 216 54 234 57
rect 258 54 276 57
rect 303 54 318 57
rect 345 54 360 57
rect 387 54 402 57
rect 429 54 450 57
rect 0 51 24 54
rect 45 51 51 54
rect 57 51 66 54
rect 87 51 96 54
rect 102 51 108 54
rect 129 51 138 54
rect 144 51 150 54
rect 171 51 180 54
rect 186 51 195 54
rect 213 51 222 54
rect 228 51 237 54
rect 255 51 264 54
rect 270 51 279 54
rect 300 51 306 54
rect 312 51 321 54
rect 342 51 348 54
rect 354 51 363 54
rect 384 51 393 54
rect 399 51 405 54
rect 426 51 450 54
rect 0 24 15 51
rect 18 48 27 51
rect 42 48 48 51
rect 60 48 69 51
rect 84 48 93 51
rect 105 48 111 51
rect 126 48 135 51
rect 147 48 153 51
rect 168 48 177 51
rect 189 48 198 51
rect 210 48 219 51
rect 231 48 240 51
rect 252 48 261 51
rect 273 48 282 51
rect 297 48 303 51
rect 315 48 324 51
rect 339 48 345 51
rect 357 48 366 51
rect 381 48 390 51
rect 402 48 408 51
rect 423 48 432 51
rect 21 45 30 48
rect 39 45 45 48
rect 63 45 72 48
rect 81 45 90 48
rect 108 45 114 48
rect 123 45 132 48
rect 150 45 156 48
rect 165 45 174 48
rect 192 45 201 48
rect 207 45 216 48
rect 234 45 243 48
rect 249 45 258 48
rect 276 45 285 48
rect 294 45 300 48
rect 318 45 327 48
rect 336 45 342 48
rect 360 45 369 48
rect 378 45 387 48
rect 405 45 411 48
rect 420 45 429 48
rect 24 42 42 45
rect 66 42 87 45
rect 111 42 129 45
rect 153 42 171 45
rect 195 42 213 45
rect 237 42 255 45
rect 279 42 297 45
rect 321 42 339 45
rect 363 42 384 45
rect 408 42 426 45
rect 27 39 39 42
rect 69 39 84 42
rect 114 39 126 42
rect 30 36 39 39
rect 72 36 81 39
rect 114 36 123 39
rect 156 36 168 42
rect 198 36 210 42
rect 240 36 252 42
rect 282 36 294 42
rect 324 39 336 42
rect 366 39 381 42
rect 411 39 423 42
rect 327 36 336 39
rect 369 36 378 39
rect 411 36 420 39
rect 27 33 42 36
rect 69 33 84 36
rect 111 33 126 36
rect 153 33 168 36
rect 195 33 213 36
rect 237 33 255 36
rect 282 33 297 36
rect 324 33 339 36
rect 366 33 381 36
rect 408 33 423 36
rect 24 30 30 33
rect 36 30 45 33
rect 66 30 75 33
rect 78 30 87 33
rect 108 30 117 33
rect 123 30 129 33
rect 150 30 159 33
rect 165 30 171 33
rect 192 30 201 33
rect 207 30 216 33
rect 234 30 243 33
rect 249 30 258 33
rect 279 30 285 33
rect 291 30 300 33
rect 321 30 327 33
rect 333 30 342 33
rect 363 30 372 33
rect 375 30 384 33
rect 405 30 414 33
rect 420 30 426 33
rect 21 27 27 30
rect 39 27 48 30
rect 63 27 72 30
rect 81 27 90 30
rect 105 27 114 30
rect 126 27 132 30
rect 147 27 156 30
rect 168 27 174 30
rect 189 27 198 30
rect 210 27 219 30
rect 231 27 240 30
rect 252 27 261 30
rect 276 27 282 30
rect 294 27 303 30
rect 318 27 324 30
rect 336 27 345 30
rect 360 27 369 30
rect 378 27 387 30
rect 402 27 411 30
rect 423 27 429 30
rect 18 24 24 27
rect 42 24 51 27
rect 60 24 69 27
rect 84 24 93 27
rect 102 24 111 27
rect 129 24 135 27
rect 144 24 153 27
rect 171 24 177 27
rect 186 24 195 27
rect 213 24 222 27
rect 228 24 237 27
rect 255 24 264 27
rect 273 24 279 27
rect 297 24 306 27
rect 315 24 321 27
rect 339 24 348 27
rect 357 24 366 27
rect 381 24 390 27
rect 399 24 408 27
rect 426 24 432 27
rect 435 24 450 51
rect 0 21 21 24
rect 45 21 66 24
rect 87 21 108 24
rect 132 21 150 24
rect 174 21 180 24
rect 183 21 192 24
rect 216 21 234 24
rect 258 21 267 24
rect 270 21 276 24
rect 300 21 309 24
rect 312 21 318 24
rect 342 21 363 24
rect 384 21 405 24
rect 429 21 450 24
rect 0 18 18 21
rect 48 18 63 21
rect 90 18 105 21
rect 135 18 147 21
rect 177 18 189 21
rect 219 18 231 21
rect 261 18 273 21
rect 303 18 315 21
rect 345 18 360 21
rect 387 18 402 21
rect 432 18 450 21
rect 0 3 450 18
<< end >>
