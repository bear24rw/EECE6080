magic
tech scmos
timestamp 1383892845
<< metal2 >>
rect 1023 4743 1277 4997
rect 1323 4743 1577 4997
rect 1623 4743 1877 4997
rect 1923 4743 2177 4997
rect 2223 4743 2477 4997
rect 2523 4743 2777 4997
rect 2823 4743 3077 4997
rect 3123 4743 3377 4997
rect 3423 4743 3677 4997
rect 3723 4743 3977 4997
rect 3 3723 257 3977
rect 4743 3723 4997 3977
rect 3 3423 257 3677
rect 4743 3423 4997 3677
rect 3 3123 257 3377
rect 4743 3123 4997 3377
rect 3 2823 257 3077
rect 4743 2823 4997 3077
rect 3 2523 257 2777
rect 4743 2523 4997 2777
rect 3 2223 257 2477
rect 4743 2223 4997 2477
rect 3 1923 257 2177
rect 4743 1923 4997 2177
rect 3 1623 257 1877
rect 4743 1623 4997 1877
rect 3 1323 257 1577
rect 4743 1323 4997 1577
rect 3 1023 257 1277
rect 4743 1023 4997 1277
rect 1023 3 1277 257
rect 1323 3 1577 257
rect 1623 3 1877 257
rect 1923 3 2177 257
rect 2223 3 2477 257
rect 2523 3 2777 257
rect 2823 3 3077 257
rect 3123 3 3377 257
rect 3423 3 3677 257
rect 3723 3 3977 257
<< labels >>
rlabel metal2 3 1023 257 1277 0 SCLKI
rlabel metal2 3 1323 257 1577 0 LDI
rlabel metal2 3 1623 257 1877 0 SI
rlabel metal2 3 1923 257 2177 0 TESTI
rlabel metal2 3 2223 257 2477 0 PSI
rlabel metal2 3 2523 257 2777 0 PCLKI
rlabel metal2 3 2823 257 3077 0 TIO
rlabel metal2 3 3123 257 3377 0 TII
rlabel metal2 3 3423 257 3677 0 TPQI
rlabel metal2 3 3723 257 3977 0 TPCI
rlabel metal2 1023 4743 1277 4997 0 TPZI
rlabel metal2 1323 4743 1577 4997 0 TPWI
rlabel metal2 1623 4743 1877 4997 0 TPZO
rlabel metal2 1923 4743 2177 4997 0 TPQO
rlabel metal2 2223 4743 2477 4997 0 VDD
rlabel metal2 2523 4743 2777 4997 0 TSSI
rlabel metal2 2823 4743 3077 4997 0 TSLDI
rlabel metal2 3123 4743 3377 4997 0 TSCI
rlabel metal2 3423 4743 3677 4997 0 TSZ
rlabel metal2 3723 4743 3977 4997 0 TSSO
rlabel metal2 4743 3723 4997 3977 0 TFQ
rlabel metal2 4743 3423 4997 3677 0 TFD
rlabel metal2 4743 3123 4997 3377 0 TFC
rlabel metal2 4743 2823 4997 3077 0 NC
rlabel metal2 4743 2523 4997 2777 0 PCLKO
rlabel metal2 4743 2223 4997 2477 0 PSO
rlabel metal2 4743 1923 4997 2177 0 TESTO
rlabel metal2 4743 1623 4997 1877 0 SO
rlabel metal2 4743 1323 4997 1577 0 LDO
rlabel metal2 4743 1023 4997 1277 0 SCLKO
rlabel metal2 3723 3 3977 257 0 W15
rlabel metal2 3423 3 3677 257 0 W14
rlabel metal2 3123 3 3377 257 0 W13
rlabel metal2 2823 3 3077 257 0 W12
rlabel metal2 2523 3 2777 257 0 GND
rlabel metal2 2223 3 2477 257 0 W4
rlabel metal2 1923 3 2177 257 0 W3
rlabel metal2 1623 3 1877 257 0 W2
rlabel metal2 1323 3 1577 257 0 W1
rlabel metal2 1023 3 1277 257 0 W0
<< end >>
