magic
tech scmos
timestamp 1383914834
<< metal1 >>
rect 20 236 1920 272
rect 20 88 268 236
rect 304 232 352 236
rect 304 228 348 232
rect 304 224 344 228
rect 304 220 340 224
rect 304 212 336 220
rect 304 208 332 212
rect 304 204 328 208
rect 304 88 324 204
rect 416 200 436 236
rect 528 200 548 236
rect 612 232 692 236
rect 752 232 800 236
rect 616 228 688 232
rect 752 228 796 232
rect 624 224 684 228
rect 628 220 684 224
rect 752 224 792 228
rect 752 220 788 224
rect 632 216 680 220
rect 636 212 676 216
rect 640 208 676 212
rect 752 212 784 220
rect 752 208 780 212
rect 640 204 672 208
rect 752 204 776 208
rect 364 88 380 200
rect 416 88 464 200
rect 20 68 464 88
rect 500 88 548 200
rect 588 176 604 200
rect 640 196 668 204
rect 712 196 716 204
rect 640 192 664 196
rect 708 192 716 196
rect 640 160 660 192
rect 704 184 716 192
rect 700 176 716 184
rect 632 152 660 160
rect 588 144 592 148
rect 636 144 660 152
rect 588 140 596 144
rect 588 136 600 140
rect 588 88 604 136
rect 500 68 604 88
rect 640 88 660 144
rect 700 88 716 152
rect 752 88 772 204
rect 812 88 828 200
rect 864 88 884 236
rect 976 200 996 236
rect 924 176 996 200
rect 1036 176 1052 236
rect 1088 200 1308 236
rect 1372 232 1448 236
rect 1376 228 1444 232
rect 1376 224 1440 228
rect 1380 220 1440 224
rect 1384 216 1436 220
rect 1384 212 1432 216
rect 1388 208 1428 212
rect 1392 204 1424 208
rect 1392 200 1420 204
rect 1088 184 1368 200
rect 1396 192 1420 200
rect 1088 180 1180 184
rect 1084 176 1180 180
rect 944 152 996 176
rect 1080 172 1180 176
rect 1076 168 1180 172
rect 1072 160 1180 168
rect 1068 156 1180 160
rect 924 148 1020 152
rect 1088 148 1180 156
rect 1216 176 1368 184
rect 1216 148 1308 176
rect 1400 148 1420 192
rect 924 144 1016 148
rect 924 140 1012 144
rect 924 136 1008 140
rect 924 132 1004 136
rect 924 128 1000 132
rect 924 124 996 128
rect 976 88 996 124
rect 1036 88 1052 132
rect 1088 88 1308 148
rect 1340 120 1420 148
rect 1460 120 1476 200
rect 1400 88 1420 120
rect 1512 116 1532 236
rect 1508 112 1532 116
rect 1504 108 1532 112
rect 1500 104 1532 108
rect 1496 100 1532 104
rect 1492 96 1532 100
rect 1488 92 1532 96
rect 1484 88 1532 92
rect 1568 200 1588 236
rect 1652 232 1920 236
rect 1656 224 1920 232
rect 1660 220 1920 224
rect 1664 212 1920 220
rect 1668 208 1920 212
rect 1672 200 1920 208
rect 1568 176 1644 200
rect 1676 192 1920 200
rect 1568 148 1624 176
rect 1568 120 1644 148
rect 1568 88 1588 120
rect 1680 108 1920 192
rect 1676 104 1920 108
rect 1672 100 1920 104
rect 1668 96 1920 100
rect 1664 92 1920 96
rect 1660 88 1920 92
rect 640 68 1920 88
rect 20 24 1920 68
<< metal2 >>
rect 0 272 1940 292
rect 0 268 32 272
rect 48 268 64 272
rect 72 268 88 272
rect 104 268 120 272
rect 128 268 144 272
rect 160 268 176 272
rect 184 268 200 272
rect 216 268 232 272
rect 240 268 256 272
rect 272 268 288 272
rect 296 268 312 272
rect 328 268 348 272
rect 352 268 368 272
rect 388 268 404 272
rect 408 268 428 272
rect 444 268 460 272
rect 468 268 484 272
rect 500 268 516 272
rect 524 268 540 272
rect 556 268 572 272
rect 580 268 596 272
rect 612 268 628 272
rect 636 268 652 272
rect 668 268 684 272
rect 692 268 708 272
rect 724 268 744 272
rect 748 268 764 272
rect 784 268 800 272
rect 804 268 824 272
rect 840 268 856 272
rect 864 268 880 272
rect 896 268 912 272
rect 920 268 936 272
rect 952 268 968 272
rect 976 268 992 272
rect 1008 268 1024 272
rect 1032 268 1048 272
rect 1064 268 1080 272
rect 1088 268 1104 272
rect 1120 268 1140 272
rect 1144 268 1160 272
rect 1180 268 1196 272
rect 1200 268 1220 272
rect 1236 268 1252 272
rect 1260 268 1276 272
rect 1292 268 1308 272
rect 1316 268 1332 272
rect 1348 268 1364 272
rect 1372 268 1388 272
rect 1404 268 1420 272
rect 1428 268 1444 272
rect 1460 268 1476 272
rect 1484 268 1500 272
rect 1516 268 1536 272
rect 1540 268 1556 272
rect 1576 268 1592 272
rect 1596 268 1616 272
rect 1632 268 1648 272
rect 1656 268 1672 272
rect 1688 268 1704 272
rect 1712 268 1728 272
rect 1744 268 1760 272
rect 1768 268 1784 272
rect 1800 268 1816 272
rect 1824 268 1840 272
rect 1856 268 1872 272
rect 1880 268 1896 272
rect 1912 268 1940 272
rect 0 264 28 268
rect 52 264 84 268
rect 108 264 140 268
rect 164 264 196 268
rect 220 264 252 268
rect 276 264 308 268
rect 332 264 364 268
rect 392 264 424 268
rect 448 264 480 268
rect 504 264 536 268
rect 560 264 592 268
rect 616 264 648 268
rect 672 264 704 268
rect 728 264 760 268
rect 788 264 820 268
rect 844 264 876 268
rect 900 264 932 268
rect 956 264 988 268
rect 1012 264 1044 268
rect 1068 264 1100 268
rect 1124 264 1156 268
rect 1184 264 1216 268
rect 1240 264 1272 268
rect 1296 264 1328 268
rect 1352 264 1384 268
rect 1408 264 1440 268
rect 1464 264 1496 268
rect 1520 264 1552 268
rect 1580 264 1612 268
rect 1636 264 1668 268
rect 1692 264 1724 268
rect 1748 264 1780 268
rect 1804 264 1836 268
rect 1860 264 1892 268
rect 1916 264 1940 268
rect 0 260 24 264
rect 56 260 80 264
rect 112 260 136 264
rect 168 260 192 264
rect 224 260 248 264
rect 280 260 304 264
rect 336 260 360 264
rect 0 256 20 260
rect 56 256 76 260
rect 112 256 132 260
rect 172 256 192 260
rect 228 256 248 260
rect 284 256 304 260
rect 340 256 360 260
rect 396 260 420 264
rect 452 260 476 264
rect 508 260 532 264
rect 564 260 588 264
rect 620 260 644 264
rect 676 260 700 264
rect 732 260 756 264
rect 396 256 416 260
rect 452 256 472 260
rect 508 256 528 260
rect 568 256 588 260
rect 624 256 644 260
rect 680 256 700 260
rect 736 256 756 260
rect 792 260 816 264
rect 848 260 872 264
rect 904 260 928 264
rect 960 260 984 264
rect 1016 260 1040 264
rect 1072 260 1096 264
rect 1128 260 1152 264
rect 792 256 812 260
rect 848 256 868 260
rect 904 256 924 260
rect 964 256 980 260
rect 1020 256 1040 260
rect 1076 256 1096 260
rect 1132 256 1152 260
rect 1188 260 1212 264
rect 1244 260 1268 264
rect 1300 260 1324 264
rect 1356 260 1380 264
rect 1412 260 1436 264
rect 1468 260 1492 264
rect 1524 260 1548 264
rect 1188 256 1208 260
rect 1244 256 1264 260
rect 1300 256 1320 260
rect 1356 256 1376 260
rect 1416 256 1436 260
rect 1472 256 1492 260
rect 1528 256 1548 260
rect 1584 260 1608 264
rect 1640 260 1664 264
rect 1696 260 1720 264
rect 1752 260 1776 264
rect 1808 260 1832 264
rect 1864 260 1888 264
rect 1584 256 1604 260
rect 1640 256 1660 260
rect 1696 256 1716 260
rect 1752 256 1772 260
rect 1812 256 1832 260
rect 1868 256 1888 260
rect 0 252 24 256
rect 56 252 80 256
rect 112 252 136 256
rect 168 252 192 256
rect 224 252 248 256
rect 280 252 304 256
rect 336 252 364 256
rect 392 252 420 256
rect 452 252 476 256
rect 508 252 532 256
rect 564 252 588 256
rect 620 252 644 256
rect 676 252 700 256
rect 732 252 760 256
rect 788 252 816 256
rect 848 252 872 256
rect 904 252 928 256
rect 960 252 984 256
rect 1016 252 1040 256
rect 1072 252 1096 256
rect 1128 252 1156 256
rect 1184 252 1212 256
rect 1244 252 1268 256
rect 1300 252 1324 256
rect 1356 252 1380 256
rect 1412 252 1436 256
rect 1468 252 1492 256
rect 1524 252 1552 256
rect 1580 252 1608 256
rect 1640 252 1664 256
rect 1696 252 1720 256
rect 1752 252 1776 256
rect 1808 252 1832 256
rect 1864 252 1888 256
rect 1920 252 1940 264
rect 0 248 28 252
rect 52 248 84 252
rect 108 248 140 252
rect 164 248 196 252
rect 220 248 252 252
rect 276 248 308 252
rect 332 248 368 252
rect 388 248 424 252
rect 448 248 480 252
rect 504 248 536 252
rect 560 248 592 252
rect 616 248 648 252
rect 672 248 704 252
rect 728 248 764 252
rect 784 248 820 252
rect 844 248 876 252
rect 900 248 932 252
rect 956 248 988 252
rect 1012 248 1044 252
rect 1068 248 1100 252
rect 1124 248 1160 252
rect 1180 248 1216 252
rect 1240 248 1272 252
rect 1296 248 1328 252
rect 1352 248 1384 252
rect 1408 248 1440 252
rect 1464 248 1496 252
rect 1520 248 1556 252
rect 1576 248 1612 252
rect 1636 248 1668 252
rect 1692 248 1724 252
rect 1748 248 1780 252
rect 1804 248 1836 252
rect 1860 248 1892 252
rect 1916 248 1940 252
rect 0 244 32 248
rect 48 244 64 248
rect 72 244 88 248
rect 104 244 120 248
rect 128 244 144 248
rect 160 244 176 248
rect 184 244 200 248
rect 216 244 232 248
rect 240 244 256 248
rect 272 244 288 248
rect 296 244 312 248
rect 328 244 344 248
rect 352 244 372 248
rect 384 244 404 248
rect 412 244 428 248
rect 444 244 460 248
rect 468 244 484 248
rect 500 244 516 248
rect 524 244 540 248
rect 556 244 572 248
rect 580 244 596 248
rect 612 244 628 248
rect 636 244 652 248
rect 668 247 684 248
rect 668 244 681 247
rect 692 244 708 248
rect 724 244 740 248
rect 748 244 768 248
rect 780 244 800 248
rect 808 244 824 248
rect 840 244 856 248
rect 864 244 880 248
rect 896 244 912 248
rect 920 244 936 248
rect 952 244 968 248
rect 976 244 992 248
rect 1008 244 1024 248
rect 1032 244 1048 248
rect 1064 244 1080 248
rect 1088 244 1104 248
rect 1120 244 1136 248
rect 1144 244 1164 248
rect 1176 244 1196 248
rect 1204 244 1220 248
rect 1236 244 1252 248
rect 1260 244 1276 248
rect 1292 244 1308 248
rect 1316 244 1332 248
rect 1348 244 1364 248
rect 1372 244 1388 248
rect 1404 244 1420 248
rect 1428 244 1444 248
rect 1460 244 1476 248
rect 1484 244 1500 248
rect 1516 244 1532 248
rect 1540 244 1560 248
rect 1572 244 1592 248
rect 1600 244 1616 248
rect 1632 244 1648 248
rect 1656 244 1672 248
rect 1688 244 1704 248
rect 1712 244 1728 248
rect 1744 244 1760 248
rect 1768 244 1784 248
rect 1800 244 1816 248
rect 1824 244 1840 248
rect 1856 244 1872 248
rect 1880 244 1896 248
rect 1912 244 1940 248
rect 0 240 36 244
rect 44 240 60 244
rect 76 240 92 244
rect 100 240 116 244
rect 132 240 148 244
rect 156 240 172 244
rect 188 240 204 244
rect 212 240 228 244
rect 244 240 316 244
rect 324 240 340 244
rect 348 240 624 244
rect 640 240 656 244
rect 664 243 680 244
rect 664 240 677 243
rect 684 240 772 244
rect 776 240 1108 244
rect 1116 240 1132 244
rect 1148 240 1168 244
rect 1172 240 1192 244
rect 1208 240 1224 244
rect 1232 240 1248 244
rect 1264 240 1280 244
rect 1288 240 1392 244
rect 1400 240 1416 244
rect 1432 240 1676 244
rect 1684 240 1700 244
rect 1716 240 1732 244
rect 1740 240 1756 244
rect 1772 240 1788 244
rect 1796 240 1812 244
rect 1828 240 1844 244
rect 1852 240 1868 244
rect 1884 240 1900 244
rect 1908 240 1940 244
rect 0 220 20 240
rect 24 236 56 240
rect 80 236 112 240
rect 136 236 168 240
rect 192 236 224 240
rect 248 236 336 240
rect 344 236 624 240
rect 644 236 676 240
rect 680 236 1128 240
rect 1152 236 1188 240
rect 1212 236 1244 240
rect 1268 236 1412 240
rect 1436 236 1696 240
rect 1720 236 1752 240
rect 1776 236 1808 240
rect 1832 236 1864 240
rect 1888 236 1940 240
rect 28 232 52 236
rect 84 232 108 236
rect 140 232 164 236
rect 196 232 220 236
rect 28 228 48 232
rect 84 228 104 232
rect 140 228 160 232
rect 200 228 216 232
rect 28 224 52 228
rect 84 224 108 228
rect 140 224 164 228
rect 196 224 220 228
rect 252 224 268 236
rect 24 220 56 224
rect 80 220 112 224
rect 136 220 168 224
rect 192 220 224 224
rect 248 220 268 224
rect 0 216 36 220
rect 44 216 60 220
rect 76 216 92 220
rect 100 216 116 220
rect 132 216 148 220
rect 156 216 172 220
rect 188 216 204 220
rect 212 216 228 220
rect 244 216 268 220
rect 0 212 32 216
rect 48 212 64 216
rect 72 212 88 216
rect 104 212 120 216
rect 128 212 144 216
rect 160 212 176 216
rect 184 212 200 216
rect 216 212 232 216
rect 240 212 268 216
rect 0 208 28 212
rect 52 208 84 212
rect 108 208 140 212
rect 164 208 196 212
rect 220 208 268 212
rect 0 204 24 208
rect 56 204 80 208
rect 112 204 136 208
rect 168 204 192 208
rect 224 204 248 208
rect 0 200 20 204
rect 56 200 76 204
rect 112 200 132 204
rect 172 200 192 204
rect 228 200 248 204
rect 0 196 24 200
rect 56 196 80 200
rect 112 196 136 200
rect 168 196 192 200
rect 224 196 248 200
rect 252 196 268 208
rect 0 192 28 196
rect 52 192 84 196
rect 108 192 140 196
rect 164 192 196 196
rect 220 192 268 196
rect 0 188 32 192
rect 48 188 64 192
rect 72 188 88 192
rect 104 188 120 192
rect 128 188 144 192
rect 160 188 176 192
rect 184 188 200 192
rect 216 188 232 192
rect 240 188 268 192
rect 0 184 36 188
rect 44 184 60 188
rect 76 184 92 188
rect 100 184 116 188
rect 132 184 148 188
rect 156 184 172 188
rect 188 184 204 188
rect 212 184 228 188
rect 244 184 268 188
rect 0 180 56 184
rect 80 180 112 184
rect 136 180 168 184
rect 192 180 224 184
rect 248 180 268 184
rect 0 164 20 180
rect 24 176 52 180
rect 84 176 108 180
rect 140 176 164 180
rect 196 176 220 180
rect 28 172 48 176
rect 84 172 104 176
rect 140 172 160 176
rect 200 172 220 176
rect 28 168 52 172
rect 84 168 108 172
rect 140 168 164 172
rect 196 168 220 172
rect 252 168 268 180
rect 24 164 56 168
rect 80 164 112 168
rect 136 164 168 168
rect 192 164 224 168
rect 248 164 268 168
rect 0 160 36 164
rect 40 160 60 164
rect 76 160 92 164
rect 100 160 116 164
rect 132 160 148 164
rect 156 160 172 164
rect 188 160 204 164
rect 212 160 228 164
rect 244 160 268 164
rect 0 156 32 160
rect 44 156 64 160
rect 72 156 88 160
rect 104 156 120 160
rect 128 156 144 160
rect 160 156 176 160
rect 184 156 200 160
rect 216 156 232 160
rect 240 156 268 160
rect 0 152 28 156
rect 48 152 84 156
rect 108 152 140 156
rect 164 152 196 156
rect 220 152 268 156
rect 0 148 24 152
rect 52 148 80 152
rect 112 148 136 152
rect 0 140 20 148
rect 56 144 76 148
rect 112 144 132 148
rect 56 140 80 144
rect 112 140 136 144
rect 168 140 192 152
rect 224 148 248 152
rect 228 144 248 148
rect 224 140 248 144
rect 252 140 268 152
rect 0 136 24 140
rect 52 136 84 140
rect 108 136 140 140
rect 164 136 196 140
rect 220 136 268 140
rect 0 132 28 136
rect 48 132 64 136
rect 68 132 88 136
rect 104 132 120 136
rect 128 132 144 136
rect 160 132 176 136
rect 184 132 200 136
rect 216 132 232 136
rect 240 132 268 136
rect 0 128 32 132
rect 44 128 60 132
rect 72 128 92 132
rect 100 128 116 132
rect 132 128 148 132
rect 156 128 172 132
rect 188 128 204 132
rect 212 128 228 132
rect 244 128 268 132
rect 0 124 56 128
rect 76 124 112 128
rect 136 124 168 128
rect 192 124 224 128
rect 248 124 268 128
rect 0 108 20 124
rect 24 120 52 124
rect 80 120 108 124
rect 140 120 164 124
rect 196 120 220 124
rect 28 112 48 120
rect 84 116 104 120
rect 140 116 160 120
rect 200 116 220 120
rect 84 112 108 116
rect 140 112 164 116
rect 196 112 220 116
rect 252 112 268 124
rect 24 108 52 112
rect 80 108 112 112
rect 136 108 168 112
rect 192 108 224 112
rect 248 108 268 112
rect 0 104 36 108
rect 40 104 56 108
rect 76 104 92 108
rect 96 104 116 108
rect 132 104 148 108
rect 156 104 172 108
rect 188 104 204 108
rect 212 104 228 108
rect 244 104 268 108
rect 0 100 32 104
rect 44 100 60 104
rect 72 100 88 104
rect 100 100 120 104
rect 128 100 144 104
rect 160 100 176 104
rect 184 100 200 104
rect 216 100 232 104
rect 240 100 268 104
rect 0 96 28 100
rect 48 96 84 100
rect 104 96 140 100
rect 164 96 196 100
rect 220 96 268 100
rect 0 92 24 96
rect 52 92 80 96
rect 108 92 136 96
rect 0 84 20 92
rect 56 84 76 92
rect 112 88 132 92
rect 112 84 136 88
rect 168 84 192 96
rect 224 92 268 96
rect 228 88 248 92
rect 224 84 248 88
rect 252 88 268 92
rect 304 228 332 236
rect 340 232 352 236
rect 336 228 348 232
rect 304 224 344 228
rect 304 220 340 224
rect 304 212 316 220
rect 324 216 336 220
rect 320 212 336 216
rect 304 208 328 212
rect 304 88 324 208
rect 416 200 436 236
rect 528 200 548 236
rect 612 232 628 236
rect 648 232 672 236
rect 680 232 688 236
rect 752 232 800 236
rect 620 228 632 232
rect 652 228 672 232
rect 676 228 684 232
rect 624 224 636 228
rect 648 224 684 228
rect 752 228 796 232
rect 752 224 792 228
rect 628 220 680 224
rect 636 216 656 220
rect 664 216 680 220
rect 752 220 788 224
rect 636 212 652 216
rect 364 88 380 200
rect 416 164 464 200
rect 416 160 432 164
rect 436 160 464 164
rect 416 128 428 160
rect 440 156 464 160
rect 444 152 464 156
rect 448 136 464 152
rect 444 132 464 136
rect 440 128 464 132
rect 416 120 464 128
rect 416 112 444 120
rect 448 112 464 120
rect 416 108 464 112
rect 416 104 432 108
rect 436 104 464 108
rect 416 88 428 104
rect 440 100 464 104
rect 444 96 464 100
rect 252 84 428 88
rect 0 80 24 84
rect 52 80 80 84
rect 108 80 140 84
rect 164 80 196 84
rect 220 80 428 84
rect 448 80 464 96
rect 0 76 28 80
rect 48 76 64 80
rect 68 76 84 80
rect 104 76 120 80
rect 124 76 144 80
rect 160 76 200 80
rect 216 76 236 80
rect 240 76 428 80
rect 444 76 464 80
rect 0 72 32 76
rect 44 72 60 76
rect 72 72 88 76
rect 100 72 116 76
rect 128 72 148 76
rect 156 72 172 76
rect 188 72 204 76
rect 212 72 232 76
rect 244 72 428 76
rect 440 72 464 76
rect 0 68 56 72
rect 76 68 112 72
rect 132 68 168 72
rect 192 68 228 72
rect 248 68 464 72
rect 500 172 548 200
rect 588 176 604 200
rect 640 196 652 212
rect 664 208 676 216
rect 752 212 784 220
rect 752 208 776 212
rect 660 204 672 208
rect 656 200 668 204
rect 656 196 664 200
rect 712 196 716 200
rect 640 192 664 196
rect 708 192 716 196
rect 500 160 512 172
rect 532 164 548 172
rect 528 160 548 164
rect 640 160 660 192
rect 704 184 716 192
rect 700 176 716 184
rect 500 156 516 160
rect 524 156 548 160
rect 500 148 548 156
rect 632 152 660 160
rect 500 144 528 148
rect 532 144 548 148
rect 636 144 660 152
rect 500 136 548 144
rect 500 132 516 136
rect 524 132 548 136
rect 500 104 512 132
rect 528 128 548 132
rect 532 108 548 128
rect 528 104 548 108
rect 500 100 516 104
rect 524 100 548 104
rect 500 92 548 100
rect 500 88 528 92
rect 532 88 548 92
rect 588 140 592 144
rect 588 136 596 140
rect 588 132 600 136
rect 588 88 604 132
rect 500 80 604 88
rect 500 76 516 80
rect 520 76 604 80
rect 500 68 512 76
rect 524 72 604 76
rect 528 68 604 72
rect 640 88 660 144
rect 700 148 704 152
rect 700 88 716 148
rect 752 88 772 208
rect 812 88 828 200
rect 864 88 884 236
rect 976 200 996 236
rect 924 176 996 200
rect 1036 176 1052 236
rect 1088 232 1124 236
rect 1156 232 1184 236
rect 1216 232 1240 236
rect 1088 228 1100 232
rect 1104 228 1124 232
rect 1160 228 1180 232
rect 1216 228 1236 232
rect 1088 224 1124 228
rect 1156 224 1184 228
rect 1216 224 1240 228
rect 1272 224 1308 236
rect 1376 228 1408 236
rect 1436 232 1448 236
rect 1432 228 1444 232
rect 1088 220 1128 224
rect 1152 220 1188 224
rect 1212 220 1244 224
rect 1268 220 1308 224
rect 1380 224 1408 228
rect 1428 224 1440 228
rect 1380 220 1412 224
rect 1424 220 1440 224
rect 1088 216 1108 220
rect 1116 216 1132 220
rect 1148 216 1168 220
rect 1172 216 1192 220
rect 1208 216 1224 220
rect 1232 216 1248 220
rect 1264 216 1280 220
rect 1288 216 1308 220
rect 1088 212 1104 216
rect 1120 212 1136 216
rect 1144 212 1164 216
rect 1176 212 1196 216
rect 1204 212 1220 216
rect 1236 212 1252 216
rect 1260 212 1276 216
rect 1088 192 1100 212
rect 1124 208 1160 212
rect 1180 208 1216 212
rect 1240 208 1272 212
rect 1128 204 1156 208
rect 1184 204 1212 208
rect 1244 204 1268 208
rect 1132 200 1152 204
rect 1128 196 1152 200
rect 1188 200 1208 204
rect 1244 200 1264 204
rect 1292 200 1308 216
rect 1384 212 1396 220
rect 1400 216 1416 220
rect 1420 216 1436 220
rect 1404 212 1432 216
rect 1388 208 1400 212
rect 1392 204 1400 208
rect 1408 208 1428 212
rect 1408 204 1424 208
rect 1188 196 1212 200
rect 1244 196 1268 200
rect 1124 192 1156 196
rect 1184 192 1216 196
rect 1240 192 1272 196
rect 1292 192 1368 200
rect 1396 196 1420 204
rect 1088 188 1104 192
rect 1120 188 1140 192
rect 1144 188 1160 192
rect 1168 188 1228 192
rect 1236 188 1252 192
rect 1260 188 1276 192
rect 1292 188 1364 192
rect 1088 184 1108 188
rect 1116 184 1136 188
rect 1148 184 1228 188
rect 1232 184 1248 188
rect 1264 184 1280 188
rect 1288 184 1364 188
rect 1088 180 1132 184
rect 1152 180 1180 184
rect 1084 176 1128 180
rect 1156 176 1180 180
rect 944 172 996 176
rect 1084 172 1100 176
rect 1104 172 1124 176
rect 944 168 956 172
rect 944 164 960 168
rect 944 160 964 164
rect 980 160 996 172
rect 1080 168 1124 172
rect 1160 168 1180 176
rect 1076 164 1128 168
rect 1156 164 1180 168
rect 1072 160 1112 164
rect 1116 160 1132 164
rect 1152 160 1180 164
rect 944 156 968 160
rect 976 156 996 160
rect 1068 156 1108 160
rect 1120 156 1136 160
rect 1148 156 1180 160
rect 944 152 996 156
rect 1088 152 1104 156
rect 1124 152 1160 156
rect 924 140 956 152
rect 960 148 996 152
rect 1012 148 1020 152
rect 960 144 1016 148
rect 960 140 1012 144
rect 924 136 1008 140
rect 1088 136 1100 152
rect 1128 148 1156 152
rect 1164 148 1180 156
rect 1216 180 1244 184
rect 1268 180 1364 184
rect 1216 176 1240 180
rect 1272 176 1364 180
rect 1216 172 1236 176
rect 1216 168 1240 172
rect 1272 168 1308 176
rect 1216 164 1244 168
rect 1268 164 1308 168
rect 1216 160 1248 164
rect 1264 160 1280 164
rect 1288 160 1308 164
rect 1216 148 1228 160
rect 1232 156 1252 160
rect 1260 156 1276 160
rect 1236 152 1272 156
rect 1240 148 1268 152
rect 1132 140 1152 148
rect 1128 136 1156 140
rect 924 132 968 136
rect 976 132 1004 136
rect 1088 132 1104 136
rect 1124 132 1140 136
rect 1144 132 1160 136
rect 1164 132 1228 148
rect 1244 144 1264 148
rect 1244 140 1268 144
rect 1240 136 1272 140
rect 1236 132 1252 136
rect 1256 132 1276 136
rect 1292 132 1308 160
rect 1400 148 1420 196
rect 924 128 1000 132
rect 924 124 996 128
rect 976 88 996 124
rect 1036 88 1052 132
rect 1088 128 1108 132
rect 1120 128 1136 132
rect 1148 128 1224 132
rect 1232 128 1248 132
rect 1260 128 1280 132
rect 1288 128 1308 132
rect 1344 128 1420 148
rect 1088 124 1132 128
rect 1152 124 1244 128
rect 1264 124 1308 128
rect 1088 120 1128 124
rect 1156 120 1240 124
rect 1268 120 1308 124
rect 1340 120 1420 128
rect 1460 124 1476 200
rect 1460 120 1468 124
rect 1088 112 1100 120
rect 1104 112 1124 120
rect 1160 112 1180 120
rect 1216 112 1236 120
rect 1272 112 1308 120
rect 1088 108 1128 112
rect 1156 108 1184 112
rect 1212 108 1240 112
rect 1268 108 1308 112
rect 1088 104 1112 108
rect 1116 104 1132 108
rect 1152 104 1168 108
rect 1172 104 1188 108
rect 1208 104 1224 108
rect 1228 104 1244 108
rect 1264 104 1280 108
rect 1284 104 1308 108
rect 1088 100 1108 104
rect 1120 100 1136 104
rect 1148 100 1164 104
rect 1176 100 1192 104
rect 1204 100 1220 104
rect 1232 100 1248 104
rect 1260 100 1276 104
rect 1288 100 1308 104
rect 1088 96 1104 100
rect 1124 96 1160 100
rect 1180 96 1216 100
rect 1236 96 1272 100
rect 1088 88 1100 96
rect 1128 92 1156 96
rect 1184 92 1212 96
rect 1240 92 1268 96
rect 640 80 1100 88
rect 1132 84 1152 92
rect 1188 84 1208 92
rect 1244 84 1264 92
rect 1292 88 1308 100
rect 1400 88 1420 120
rect 1512 116 1532 236
rect 1508 112 1532 116
rect 1504 108 1532 112
rect 1500 104 1532 108
rect 1496 100 1532 104
rect 1492 96 1532 100
rect 1488 92 1532 96
rect 1484 88 1512 92
rect 1516 88 1532 92
rect 1568 200 1588 236
rect 1656 232 1664 236
rect 1668 232 1692 236
rect 1724 232 1748 236
rect 1780 232 1804 236
rect 1836 232 1860 236
rect 1892 232 1916 236
rect 1656 228 1688 232
rect 1724 228 1744 232
rect 1784 228 1804 232
rect 1840 228 1860 232
rect 1896 228 1916 232
rect 1660 224 1692 228
rect 1724 224 1748 228
rect 1780 224 1804 228
rect 1836 224 1860 228
rect 1892 224 1916 228
rect 1920 224 1940 236
rect 1660 220 1696 224
rect 1720 220 1752 224
rect 1776 220 1808 224
rect 1832 220 1864 224
rect 1888 220 1940 224
rect 1664 212 1676 220
rect 1684 216 1700 220
rect 1716 216 1732 220
rect 1740 216 1756 220
rect 1772 216 1788 220
rect 1796 216 1812 220
rect 1828 216 1844 220
rect 1852 216 1868 220
rect 1884 216 1900 220
rect 1908 216 1940 220
rect 1688 212 1704 216
rect 1712 212 1728 216
rect 1744 212 1760 216
rect 1768 212 1784 216
rect 1800 212 1816 216
rect 1824 212 1840 216
rect 1856 212 1872 216
rect 1880 212 1896 216
rect 1912 212 1940 216
rect 1668 208 1680 212
rect 1692 208 1724 212
rect 1748 208 1780 212
rect 1804 208 1836 212
rect 1860 208 1892 212
rect 1916 208 1940 212
rect 1672 204 1680 208
rect 1696 204 1720 208
rect 1752 204 1776 208
rect 1808 204 1832 208
rect 1864 204 1888 208
rect 1676 200 1684 204
rect 1696 200 1716 204
rect 1752 200 1772 204
rect 1812 200 1832 204
rect 1868 200 1888 204
rect 1568 176 1644 200
rect 1676 196 1688 200
rect 1696 196 1720 200
rect 1752 196 1776 200
rect 1808 196 1832 200
rect 1864 196 1888 200
rect 1920 196 1940 208
rect 1680 192 1688 196
rect 1692 192 1724 196
rect 1748 192 1780 196
rect 1804 192 1836 196
rect 1860 192 1892 196
rect 1916 192 1940 196
rect 1680 188 1704 192
rect 1712 188 1728 192
rect 1744 188 1760 192
rect 1768 188 1784 192
rect 1800 188 1816 192
rect 1824 188 1840 192
rect 1856 188 1872 192
rect 1880 188 1896 192
rect 1912 188 1940 192
rect 1680 184 1700 188
rect 1716 184 1732 188
rect 1740 184 1756 188
rect 1772 184 1788 188
rect 1796 184 1812 188
rect 1828 184 1844 188
rect 1852 184 1868 188
rect 1884 184 1900 188
rect 1908 184 1940 188
rect 1680 180 1696 184
rect 1720 180 1752 184
rect 1776 180 1808 184
rect 1832 180 1864 184
rect 1888 180 1940 184
rect 1568 172 1624 176
rect 1568 164 1580 172
rect 1612 168 1624 172
rect 1608 164 1624 168
rect 1568 160 1584 164
rect 1604 160 1624 164
rect 1568 156 1588 160
rect 1600 156 1624 160
rect 1568 148 1624 156
rect 1680 168 1692 180
rect 1724 176 1748 180
rect 1780 176 1804 180
rect 1836 176 1860 180
rect 1892 176 1940 180
rect 1724 172 1744 176
rect 1784 172 1804 176
rect 1840 172 1860 176
rect 1896 172 1916 176
rect 1724 168 1748 172
rect 1780 168 1804 172
rect 1836 168 1860 172
rect 1892 168 1916 172
rect 1920 168 1940 176
rect 1680 164 1696 168
rect 1720 164 1752 168
rect 1776 164 1808 168
rect 1832 164 1864 168
rect 1888 164 1940 168
rect 1680 160 1700 164
rect 1716 160 1732 164
rect 1740 160 1756 164
rect 1772 160 1788 164
rect 1796 160 1812 164
rect 1828 160 1844 164
rect 1852 160 1868 164
rect 1884 160 1904 164
rect 1908 160 1940 164
rect 1680 156 1704 160
rect 1712 156 1728 160
rect 1744 156 1760 160
rect 1768 156 1784 160
rect 1800 156 1816 160
rect 1824 156 1840 160
rect 1856 156 1872 160
rect 1880 156 1900 160
rect 1912 156 1940 160
rect 1680 152 1724 156
rect 1748 152 1780 156
rect 1804 152 1836 156
rect 1860 152 1896 156
rect 1916 152 1940 156
rect 1568 140 1580 148
rect 1584 140 1604 148
rect 1608 140 1644 148
rect 1568 136 1644 140
rect 1568 132 1592 136
rect 1596 132 1644 136
rect 1568 128 1588 132
rect 1600 128 1644 132
rect 1568 120 1644 128
rect 1680 140 1692 152
rect 1696 148 1720 152
rect 1696 144 1716 148
rect 1696 140 1720 144
rect 1752 140 1776 152
rect 1808 148 1832 152
rect 1864 148 1892 152
rect 1812 144 1832 148
rect 1868 144 1888 148
rect 1808 140 1832 144
rect 1864 140 1888 144
rect 1680 136 1724 140
rect 1748 136 1780 140
rect 1804 136 1836 140
rect 1860 136 1892 140
rect 1920 136 1940 152
rect 1680 132 1704 136
rect 1712 132 1728 136
rect 1744 132 1760 136
rect 1768 132 1784 136
rect 1800 132 1816 136
rect 1824 132 1840 136
rect 1856 132 1876 136
rect 1880 132 1896 136
rect 1916 132 1940 136
rect 1680 128 1700 132
rect 1716 128 1732 132
rect 1740 128 1756 132
rect 1772 128 1788 132
rect 1796 128 1812 132
rect 1828 128 1844 132
rect 1852 128 1872 132
rect 1884 128 1900 132
rect 1912 128 1940 132
rect 1680 124 1696 128
rect 1720 124 1752 128
rect 1776 124 1808 128
rect 1832 124 1868 128
rect 1888 124 1940 128
rect 1568 88 1588 120
rect 1680 112 1692 124
rect 1724 120 1748 124
rect 1780 120 1804 124
rect 1836 120 1864 124
rect 1892 120 1940 124
rect 1724 116 1744 120
rect 1784 116 1804 120
rect 1840 116 1860 120
rect 1724 112 1748 116
rect 1780 112 1804 116
rect 1836 112 1860 116
rect 1896 112 1916 120
rect 1920 112 1940 120
rect 1680 108 1696 112
rect 1720 108 1752 112
rect 1776 108 1808 112
rect 1832 108 1864 112
rect 1892 108 1940 112
rect 1676 104 1700 108
rect 1716 104 1732 108
rect 1740 104 1756 108
rect 1772 104 1788 108
rect 1796 104 1812 108
rect 1828 104 1848 108
rect 1852 104 1868 108
rect 1888 104 1904 108
rect 1908 104 1940 108
rect 1672 100 1704 104
rect 1712 100 1728 104
rect 1744 100 1760 104
rect 1768 100 1784 104
rect 1800 100 1816 104
rect 1824 100 1844 104
rect 1856 100 1872 104
rect 1884 100 1900 104
rect 1912 100 1940 104
rect 1668 96 1724 100
rect 1748 96 1780 100
rect 1804 96 1840 100
rect 1860 96 1896 100
rect 1916 96 1940 100
rect 1664 92 1688 96
rect 1692 92 1720 96
rect 1660 88 1688 92
rect 1696 88 1716 92
rect 1292 84 1508 88
rect 1516 84 1684 88
rect 1696 84 1720 88
rect 1752 84 1776 96
rect 1808 92 1836 96
rect 1864 92 1892 96
rect 1812 88 1832 92
rect 1808 84 1832 88
rect 1868 84 1888 92
rect 1128 80 1156 84
rect 1184 80 1212 84
rect 1240 80 1268 84
rect 640 76 1104 80
rect 1124 76 1140 80
rect 1144 76 1160 80
rect 1180 76 1196 80
rect 1200 76 1216 80
rect 1236 76 1252 80
rect 1256 76 1272 80
rect 1292 76 1504 84
rect 640 72 1108 76
rect 1120 72 1136 76
rect 1148 72 1164 76
rect 1176 72 1192 76
rect 1204 72 1220 76
rect 1232 72 1248 76
rect 1260 72 1276 76
rect 1288 72 1504 76
rect 1516 80 1680 84
rect 1692 80 1724 84
rect 1748 80 1780 84
rect 1804 80 1836 84
rect 1864 80 1892 84
rect 1920 80 1940 96
rect 1516 72 1676 80
rect 1688 76 1704 80
rect 1708 76 1728 80
rect 1744 76 1784 80
rect 1800 76 1820 80
rect 1824 76 1840 80
rect 1860 76 1876 80
rect 1880 76 1896 80
rect 1916 76 1940 80
rect 1684 72 1700 76
rect 1712 72 1732 76
rect 1740 72 1756 76
rect 1772 72 1788 76
rect 1796 72 1816 76
rect 1828 72 1844 76
rect 1856 72 1872 76
rect 1884 72 1900 76
rect 1912 72 1940 76
rect 640 68 1132 72
rect 1152 68 1188 72
rect 1208 68 1244 72
rect 1264 68 1696 72
rect 1716 68 1752 72
rect 1776 68 1812 72
rect 1832 68 1868 72
rect 1888 68 1940 72
rect 0 52 20 68
rect 24 64 52 68
rect 80 64 108 68
rect 136 64 164 68
rect 196 64 224 68
rect 252 64 512 68
rect 28 56 48 64
rect 84 60 104 64
rect 140 60 160 64
rect 84 56 108 60
rect 140 56 164 60
rect 196 56 220 64
rect 252 60 444 64
rect 256 56 276 60
rect 312 56 332 60
rect 368 56 388 60
rect 424 56 444 60
rect 448 56 512 64
rect 532 60 1096 68
rect 1100 64 1128 68
rect 1156 64 1184 68
rect 1212 64 1240 68
rect 1268 64 1488 68
rect 1496 64 1692 68
rect 1720 64 1748 68
rect 536 56 560 60
rect 588 56 672 60
rect 708 56 728 60
rect 764 56 784 60
rect 820 56 840 60
rect 876 56 896 60
rect 932 56 956 60
rect 988 56 1012 60
rect 1048 56 1068 60
rect 1104 56 1124 64
rect 1160 56 1180 64
rect 1216 56 1236 64
rect 1272 60 1484 64
rect 1500 60 1664 64
rect 1272 56 1292 60
rect 1328 56 1352 60
rect 1384 56 1408 60
rect 1444 56 1464 60
rect 1500 56 1520 60
rect 1556 56 1576 60
rect 1612 56 1632 60
rect 1668 56 1688 64
rect 1724 56 1748 64
rect 1780 64 1808 68
rect 1836 64 1864 68
rect 1892 64 1940 68
rect 1780 56 1804 64
rect 1840 60 1860 64
rect 1836 56 1860 60
rect 1896 56 1916 64
rect 1920 56 1940 64
rect 24 52 52 56
rect 80 52 108 56
rect 136 52 168 56
rect 192 52 224 56
rect 252 52 280 56
rect 308 52 336 56
rect 364 52 392 56
rect 420 52 512 56
rect 532 52 564 56
rect 588 52 676 56
rect 704 52 732 56
rect 760 52 788 56
rect 816 52 844 56
rect 872 52 900 56
rect 928 52 960 56
rect 984 52 1016 56
rect 1044 52 1072 56
rect 1100 52 1128 56
rect 1156 52 1184 56
rect 1212 52 1240 56
rect 1268 52 1296 56
rect 1324 52 1356 56
rect 1380 52 1412 56
rect 1440 52 1468 56
rect 1496 52 1524 56
rect 1552 52 1580 56
rect 1608 52 1636 56
rect 1664 52 1692 56
rect 1720 52 1752 56
rect 1776 52 1808 56
rect 1836 52 1864 56
rect 1892 52 1940 56
rect 0 48 36 52
rect 40 48 56 52
rect 76 48 92 52
rect 96 48 112 52
rect 132 48 172 52
rect 188 48 228 52
rect 248 48 264 52
rect 268 48 284 52
rect 304 48 320 52
rect 324 48 340 52
rect 360 48 376 52
rect 380 48 396 52
rect 416 48 432 52
rect 436 48 512 52
rect 528 48 568 52
rect 584 48 660 52
rect 664 48 680 52
rect 700 48 716 52
rect 720 48 736 52
rect 756 48 772 52
rect 776 48 792 52
rect 812 48 828 52
rect 832 48 848 52
rect 868 48 884 52
rect 888 48 904 52
rect 924 48 964 52
rect 980 48 1020 52
rect 1040 48 1056 52
rect 1060 48 1076 52
rect 1096 48 1112 52
rect 1116 48 1132 52
rect 1152 48 1168 52
rect 1172 48 1188 52
rect 1208 48 1224 52
rect 1228 48 1244 52
rect 1264 48 1280 52
rect 1284 48 1300 52
rect 1320 48 1360 52
rect 1376 48 1416 52
rect 1436 48 1452 52
rect 1456 48 1472 52
rect 1492 48 1508 52
rect 1512 48 1528 52
rect 1548 48 1564 52
rect 1568 48 1584 52
rect 1604 48 1620 52
rect 1624 48 1640 52
rect 1660 48 1676 52
rect 1680 48 1696 52
rect 1716 48 1756 52
rect 1772 48 1812 52
rect 1832 48 1848 52
rect 1852 48 1868 52
rect 1888 48 1904 52
rect 1908 48 1940 52
rect 0 44 32 48
rect 44 44 60 48
rect 72 44 88 48
rect 100 44 116 48
rect 128 44 144 48
rect 156 44 176 48
rect 184 44 204 48
rect 216 44 232 48
rect 244 44 260 48
rect 272 44 288 48
rect 300 44 316 48
rect 328 44 344 48
rect 356 44 372 48
rect 384 44 400 48
rect 412 44 428 48
rect 440 44 512 48
rect 524 44 540 48
rect 552 44 572 48
rect 580 44 656 48
rect 668 44 684 48
rect 696 44 712 48
rect 724 44 740 48
rect 752 44 768 48
rect 780 44 796 48
rect 808 44 824 48
rect 836 44 852 48
rect 864 44 880 48
rect 892 44 908 48
rect 920 44 936 48
rect 948 44 968 48
rect 976 44 996 48
rect 1008 44 1024 48
rect 1036 44 1052 48
rect 1064 44 1080 48
rect 1092 44 1108 48
rect 1120 44 1136 48
rect 1148 44 1164 48
rect 1176 44 1192 48
rect 1204 44 1220 48
rect 1232 44 1248 48
rect 1260 44 1276 48
rect 1288 44 1304 48
rect 1316 44 1332 48
rect 1344 44 1364 48
rect 1372 44 1392 48
rect 1404 44 1420 48
rect 1432 44 1448 48
rect 1460 44 1476 48
rect 1488 44 1504 48
rect 1516 44 1532 48
rect 1544 44 1560 48
rect 1572 44 1588 48
rect 1600 44 1616 48
rect 1628 44 1644 48
rect 1656 44 1672 48
rect 1684 44 1700 48
rect 1712 44 1728 48
rect 1740 44 1760 48
rect 1768 44 1788 48
rect 1800 44 1816 48
rect 1828 44 1844 48
rect 1856 44 1872 48
rect 1884 44 1900 48
rect 1912 44 1940 48
rect 0 40 28 44
rect 48 40 84 44
rect 104 40 140 44
rect 160 40 200 44
rect 220 40 256 44
rect 276 40 312 44
rect 332 40 368 44
rect 388 40 424 44
rect 444 40 536 44
rect 556 40 652 44
rect 672 40 708 44
rect 728 40 764 44
rect 784 40 820 44
rect 840 40 876 44
rect 896 40 932 44
rect 952 40 992 44
rect 1012 40 1048 44
rect 1068 40 1104 44
rect 1124 40 1160 44
rect 1180 40 1216 44
rect 1236 40 1272 44
rect 1292 40 1328 44
rect 1348 40 1388 44
rect 1408 40 1444 44
rect 1464 40 1500 44
rect 1520 40 1556 44
rect 1576 40 1612 44
rect 1632 40 1668 44
rect 1688 40 1724 44
rect 1744 40 1784 44
rect 1804 40 1840 44
rect 1860 40 1896 44
rect 1916 40 1940 44
rect 0 36 24 40
rect 52 36 80 40
rect 108 36 136 40
rect 164 36 196 40
rect 224 36 252 40
rect 280 36 308 40
rect 336 36 364 40
rect 392 36 420 40
rect 448 36 476 40
rect 504 36 532 40
rect 560 36 592 40
rect 620 36 648 40
rect 676 36 704 40
rect 732 36 760 40
rect 788 36 816 40
rect 844 36 872 40
rect 900 36 928 40
rect 956 36 988 40
rect 1016 36 1044 40
rect 1072 36 1100 40
rect 1128 36 1156 40
rect 1184 36 1212 40
rect 1240 36 1268 40
rect 1296 36 1324 40
rect 1352 36 1384 40
rect 1412 36 1440 40
rect 1468 36 1496 40
rect 1524 36 1552 40
rect 1580 36 1608 40
rect 1636 36 1664 40
rect 1692 36 1720 40
rect 1748 36 1780 40
rect 1808 36 1836 40
rect 1864 36 1892 40
rect 0 28 20 36
rect 56 28 76 36
rect 112 28 136 36
rect 168 28 192 36
rect 224 28 248 36
rect 284 28 304 36
rect 340 28 360 36
rect 396 28 416 36
rect 452 28 472 36
rect 508 28 532 36
rect 564 28 588 36
rect 620 28 644 36
rect 680 28 700 36
rect 736 28 756 36
rect 792 28 812 36
rect 848 28 868 36
rect 904 28 928 36
rect 960 28 984 36
rect 1016 28 1040 36
rect 1076 28 1096 36
rect 1132 28 1152 36
rect 1188 28 1208 36
rect 1244 28 1264 36
rect 1300 28 1324 36
rect 1356 28 1380 36
rect 1412 28 1436 36
rect 1472 28 1492 36
rect 1528 28 1548 36
rect 1584 28 1604 36
rect 1640 28 1660 36
rect 1696 28 1720 36
rect 1752 28 1776 36
rect 1808 28 1832 36
rect 1868 28 1888 36
rect 0 24 24 28
rect 52 24 80 28
rect 108 24 136 28
rect 164 24 196 28
rect 224 24 252 28
rect 280 24 308 28
rect 336 24 364 28
rect 392 24 420 28
rect 448 24 476 28
rect 504 24 532 28
rect 560 24 592 28
rect 620 24 648 28
rect 676 24 704 28
rect 732 24 760 28
rect 788 24 816 28
rect 844 24 872 28
rect 900 24 928 28
rect 956 24 988 28
rect 1016 24 1044 28
rect 1072 24 1100 28
rect 1128 24 1156 28
rect 1184 24 1212 28
rect 1240 24 1268 28
rect 1296 24 1324 28
rect 1352 24 1384 28
rect 1412 24 1440 28
rect 1468 24 1496 28
rect 1524 24 1552 28
rect 1580 24 1608 28
rect 1636 24 1664 28
rect 1692 24 1720 28
rect 1748 24 1780 28
rect 1808 24 1836 28
rect 1864 24 1892 28
rect 1920 24 1940 40
rect 0 4 1940 24
<< end >>
