magic
tech scmos
timestamp 1383645441
<< metal1 >>
rect -4 40 3 41
<< m2contact >>
rect -141 46 -137 50
rect -133 46 -129 50
rect -109 46 -105 50
rect -83 46 -79 50
rect -75 46 -71 50
rect -51 46 -47 50
rect -1 45 3 49
rect -91 36 -87 40
rect -33 36 -29 40
<< metal2 >>
rect -145 60 -71 64
rect -145 53 -129 57
rect -133 50 -129 53
rect -125 53 -79 57
rect -141 43 -137 46
rect -125 43 -121 53
rect -83 50 -79 53
rect -141 39 -121 43
rect -125 0 -121 39
rect -75 50 -71 60
rect -25 58 -21 1674
rect 2347 1670 2445 1674
rect 2347 1636 2438 1640
rect 2347 1520 2432 1524
rect 2347 1404 2426 1408
rect 2347 1288 2420 1292
rect 2347 1172 2414 1176
rect 2347 1056 2408 1060
rect 2347 940 2402 944
rect 2347 824 2396 828
rect 2347 708 2390 712
rect 2347 592 2384 596
rect 2347 476 2378 480
rect 2347 360 2372 364
rect 2347 244 2366 248
rect 2347 128 2360 132
rect -67 54 -21 58
rect -109 0 -105 46
rect -67 40 -63 54
rect -87 36 -63 40
rect -25 46 -21 54
rect -51 0 -47 46
rect -17 45 -1 49
rect -17 40 -13 45
rect -29 36 -13 40
rect 2347 37 2354 41
rect 2350 0 2354 37
rect 2357 0 2360 128
rect 2363 0 2366 244
rect 2369 0 2372 360
rect 2375 0 2378 476
rect 2381 0 2384 592
rect 2387 0 2390 708
rect 2393 0 2396 824
rect 2399 0 2402 940
rect 2405 0 2408 1056
rect 2411 0 2414 1172
rect 2417 0 2420 1288
rect 2423 0 2426 1404
rect 2429 0 2432 1520
rect 2435 0 2438 1636
rect 2441 0 2445 1670
use mux  mux_0
timestamp 1383644076
transform 1 0 -148 0 1 0
box 0 0 73 108
use mux  mux_1
timestamp 1383644076
transform 1 0 -90 0 1 0
box 0 0 73 108
use pin_buffer  pin_buffer_0
array 0 0 46 0 14 116
timestamp 1383629942
transform 1 0 -36 0 1 0
box 0 0 46 108
use pin_row_connect  pin_row_connect_0
array 0 0 98 0 13 116
timestamp 1383629942
transform 1 0 4 0 1 0
box -8 0 2347 165
use pin_slice  pin_slice_0
array 0 14 156 0 14 116
timestamp 1383629942
transform 1 0 100 0 1 113
box -100 -113 68 -5
<< labels >>
rlabel metal2 -145 60 -141 64 0 PSI
rlabel metal2 -145 53 -141 57 0 PCLKI
<< end >>
