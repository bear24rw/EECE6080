magic
tech scmos
timestamp 1383882935
<< m2contact >>
rect -158 129 -154 133
rect -4 129 0 133
rect 150 129 154 133
rect 304 129 308 133
rect 458 129 462 133
rect 1690 129 1694 133
rect 1844 129 1848 133
rect 1998 129 2002 133
rect 2152 129 2156 133
<< metal2 >>
rect -158 133 -154 136
rect -158 42 -154 129
rect -4 133 0 136
rect -4 48 0 129
rect 150 133 154 136
rect 150 54 154 129
rect 304 133 308 136
rect 304 60 308 129
rect 458 133 462 136
rect 458 66 462 129
rect 612 72 616 136
rect 766 78 770 136
rect 920 84 924 136
rect 1074 90 1078 136
rect 1228 96 1232 136
rect 1382 102 1386 136
rect 1536 108 1540 136
rect 1690 133 1694 136
rect 1690 114 1694 129
rect 1844 133 1848 136
rect 1844 120 1848 129
rect 1998 133 2002 136
rect 2152 133 2156 136
rect 2156 129 2274 132
rect 1998 126 2002 129
rect 1998 123 2274 126
rect 1844 117 2274 120
rect 1690 111 2274 114
rect 1536 105 2274 108
rect 1382 99 2274 102
rect 1228 93 2274 96
rect 1074 87 2274 90
rect 920 81 2274 84
rect 766 75 2274 78
rect 612 69 2274 72
rect 458 63 2274 66
rect 304 57 2274 60
rect 150 51 2274 54
rect -4 45 2274 48
rect -158 39 2274 42
use mux  mux_0
timestamp 1383808422
transform 1 0 2209 0 -1 342
box 0 0 73 108
use shift_slice  shift_slice_0
array 0 15 154 0 0 108
timestamp 1383875311
transform 1 0 -181 0 1 136
box -16 0 151 108
<< end >>
